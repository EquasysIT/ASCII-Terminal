--------------------------------------------------------------
-- Engineer: A Burgess                                      --
--                                                          --
-- Design Name: Basic Computer System - WOZ ROM             --
--                                                          --
--------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity wozrom is
	port (
		clk		    : in    std_logic;
		addr		: in    std_logic_vector(8 downto 0);
		data		: out   std_logic_vector(7 downto 0)
	);
end;

architecture rtl of wozrom is
	type romdata is array(0 to 511) of std_logic_vector(7 downto 0);
	constant rom : romdata := (
		x"A0",x"7F",x"C9",x"7F",x"F0",x"18",x"C9",x"1B", -- 0x0000
		x"F0",x"03",x"C8",x"10",x"14",x"A9",x"5C",x"20", -- 0x0008
		x"FC",x"40",x"A9",x"0D",x"20",x"FC",x"40",x"A9", -- 0x0010
		x"0A",x"20",x"FC",x"40",x"A0",x"01",x"88",x"30", -- 0x0018
		x"F1",x"AD",x"E2",x"BF",x"29",x"01",x"F0",x"06", -- 0x0020
		x"AD",x"E5",x"BF",x"4C",x"38",x"40",x"AD",x"E2", -- 0x0028
		x"BF",x"29",x"02",x"F0",x"EC",x"AD",x"E6",x"BF", -- 0x0030
		x"99",x"00",x"02",x"20",x"FC",x"40",x"C9",x"0D", -- 0x0038
		x"D0",x"C0",x"A0",x"FF",x"A9",x"00",x"AA",x"0A", -- 0x0040
		x"0A",x"85",x"2B",x"C8",x"B9",x"00",x"02",x"C9", -- 0x0048
		x"0D",x"F0",x"BF",x"C9",x"2E",x"90",x"F4",x"F0", -- 0x0050
		x"EE",x"C9",x"3A",x"F0",x"EB",x"C9",x"52",x"F0", -- 0x0058
		x"3B",x"86",x"28",x"86",x"29",x"84",x"2A",x"B9", -- 0x0060
		x"00",x"02",x"49",x"30",x"C9",x"0A",x"90",x"06", -- 0x0068
		x"69",x"88",x"C9",x"FA",x"90",x"11",x"0A",x"0A", -- 0x0070
		x"0A",x"0A",x"A2",x"04",x"0A",x"26",x"28",x"26", -- 0x0078
		x"29",x"CA",x"D0",x"F8",x"C8",x"D0",x"E0",x"C4", -- 0x0080
		x"2A",x"F0",x"82",x"24",x"2B",x"50",x"10",x"A5", -- 0x0088
		x"28",x"81",x"26",x"E6",x"26",x"D0",x"B5",x"E6", -- 0x0090
		x"27",x"4C",x"4C",x"40",x"6C",x"24",x"00",x"30", -- 0x0098
		x"30",x"A2",x"02",x"B5",x"27",x"95",x"25",x"95", -- 0x00A0
		x"23",x"CA",x"D0",x"F7",x"D0",x"19",x"A9",x"0D", -- 0x00A8
		x"20",x"FC",x"40",x"A9",x"0A",x"20",x"FC",x"40", -- 0x00B0
		x"A5",x"25",x"20",x"E9",x"40",x"A5",x"24",x"20", -- 0x00B8
		x"E9",x"40",x"A9",x"3A",x"20",x"FC",x"40",x"A9", -- 0x00C0
		x"20",x"20",x"FC",x"40",x"A1",x"24",x"20",x"E9", -- 0x00C8
		x"40",x"86",x"2B",x"A5",x"24",x"C5",x"28",x"A5", -- 0x00D0
		x"25",x"E5",x"29",x"B0",x"BC",x"E6",x"24",x"D0", -- 0x00D8
		x"02",x"E6",x"25",x"A5",x"24",x"29",x"07",x"10", -- 0x00E0
		x"C3",x"48",x"4A",x"4A",x"4A",x"4A",x"20",x"F2", -- 0x00E8
		x"40",x"68",x"29",x"0F",x"09",x"30",x"C9",x"3A", -- 0x00F0
		x"90",x"02",x"69",x"06",x"48",x"AD",x"E0",x"BF", -- 0x00F8
		x"29",x"01",x"D0",x"F9",x"68",x"8D",x"E4",x"BF", -- 0x0100
		x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0108
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0110
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0118
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0120
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0128
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0130
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0138
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0140
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0148
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0150
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0158
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0160
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0168
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0170
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0178
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0180
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0188
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0190
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0198
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x01F8
	);

begin
	process(clk)
	begin
		if rising_edge(clk) then
			data <= rom(to_integer(unsigned(addr)));
		end if;
	end process;
end rtl;
