--------------------------------------------------------------
-- Engineer: A Burgess                                      --
--                                                          --
-- Design Name: Pixel Character ROM                         --
--                                                          --
-- October 2024                                             --
--------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity pixelrom is
    port (
        clk  : in  std_logic;
        addr : in  std_logic_vector(9 downto 0);
        data : out std_logic_vector(7 downto 0)
        );
end;

architecture rtl of pixelrom is

    signal rom_addr : std_logic_vector(9 downto 0);

begin

    p_addr : process(addr)
    begin
        rom_addr              <= (others => '0');
        rom_addr(9 downto 0) <= addr;
    end process;

    p_rom : process
    begin
        wait until rising_edge(clk);
        data <= (others => '0');
        case rom_addr is
            when d"0000000000" => data <= "11111111";
            when d"0000000001" => data <= "11111111";
            when d"0000000002" => data <= "11111111";
            when d"0000000003" => data <= "11111111";
            when d"0000000004" => data <= "11111111";
            when d"0000000005" => data <= "11111111";
            when d"0000000006" => data <= "11111111";
            when d"0000000007" => data <= "11111111";
            when d"0000000008" => data <= "11111111";
            when d"0000000009" => data <= "11111111";
            when d"0000000010" => data <= "11111111";
            when d"0000000011" => data <= "11111111";
            when d"0000000012" => data <= "11111111";
            when d"0000000013" => data <= "11111111";
            when d"0000000014" => data <= "11111111";
            when d"0000000015" => data <= "11111111";
            when d"0000000016" => data <= "11111111";
            when d"0000000017" => data <= "11111111";
            when d"0000000018" => data <= "11111111";
            when d"0000000019" => data <= "11111111";
            when d"0000000020" => data <= "11111111";
            when d"0000000021" => data <= "11111111";
            when d"0000000022" => data <= "11111111";
            when d"0000000023" => data <= "11111111";
            when d"0000000024" => data <= "11111111";
            when d"0000000025" => data <= "11111111";
            when d"0000000026" => data <= "11111111";
            when d"0000000027" => data <= "11111111";
            when d"0000000028" => data <= "11111111";
            when d"0000000029" => data <= "11111111";
            when d"0000000030" => data <= "11111111";
            when d"0000000031" => data <= "11111111";
            when d"0000000032" => data <= "11111111";
            when d"0000000033" => data <= "11101111";
            when d"0000000034" => data <= "11011011";
            when d"0000000035" => data <= "11011011";
            when d"0000000036" => data <= "11110111";
            when d"0000000037" => data <= "10011101";
            when d"0000000038" => data <= "11101111";
            when d"0000000039" => data <= "11110111";
            when d"0000000040" => data <= "11111011";
            when d"0000000041" => data <= "11011111";
            when d"0000000042" => data <= "11111111";
            when d"0000000043" => data <= "11111111";
            when d"0000000044" => data <= "11111111";
            when d"0000000045" => data <= "11111111";
            when d"0000000046" => data <= "11111111";
            when d"0000000047" => data <= "11111111";
            when d"0000000048" => data <= "11000011";
            when d"0000000049" => data <= "11100111";
            when d"0000000050" => data <= "11000011";
            when d"0000000051" => data <= "11000011";
            when d"0000000052" => data <= "11110111";
            when d"0000000053" => data <= "10000001";
            when d"0000000054" => data <= "11000011";
            when d"0000000055" => data <= "10000001";
            when d"0000000056" => data <= "11000011";
            when d"0000000057" => data <= "11000011";
            when d"0000000058" => data <= "11111111";
            when d"0000000059" => data <= "11111111";
            when d"0000000060" => data <= "11111111";
            when d"0000000061" => data <= "11111111";
            when d"0000000062" => data <= "11111111";
            when d"0000000063" => data <= "11000011";
            when d"0000000064" => data <= "11111111";
            when d"0000000065" => data <= "11101111";
            when d"0000000066" => data <= "11011011";
            when d"0000000067" => data <= "10000001";
            when d"0000000068" => data <= "11000001";
            when d"0000000069" => data <= "10011011";
            when d"0000000070" => data <= "11010111";
            when d"0000000071" => data <= "11101111";
            when d"0000000072" => data <= "11110111";
            when d"0000000073" => data <= "11101111";
            when d"0000000074" => data <= "11101011";
            when d"0000000075" => data <= "11110111";
            when d"0000000076" => data <= "11111111";
            when d"0000000077" => data <= "11111111";
            when d"0000000078" => data <= "11111111";
            when d"0000000079" => data <= "11111101";
            when d"0000000080" => data <= "10111001";
            when d"0000000081" => data <= "11010111";
            when d"0000000082" => data <= "10111101";
            when d"0000000083" => data <= "10111101";
            when d"0000000084" => data <= "11100111";
            when d"0000000085" => data <= "10111111";
            when d"0000000086" => data <= "10111111";
            when d"0000000087" => data <= "11111101";
            when d"0000000088" => data <= "10111101";
            when d"0000000089" => data <= "10111101";
            when d"0000000090" => data <= "11111111";
            when d"0000000091" => data <= "11101111";
            when d"0000000092" => data <= "11111011";
            when d"0000000093" => data <= "11111111";
            when d"0000000094" => data <= "11101111";
            when d"0000000095" => data <= "10111101";
            when d"0000000096" => data <= "11111111";
            when d"0000000097" => data <= "11101111";
            when d"0000000098" => data <= "11111111";
            when d"0000000099" => data <= "11011011";
            when d"0000000100" => data <= "11010111";
            when d"0000000101" => data <= "11110111";
            when d"0000000102" => data <= "11101111";
            when d"0000000103" => data <= "11111111";
            when d"0000000104" => data <= "11110111";
            when d"0000000105" => data <= "11101111";
            when d"0000000106" => data <= "11110111";
            when d"0000000107" => data <= "11110111";
            when d"0000000108" => data <= "11111111";
            when d"0000000109" => data <= "11111111";
            when d"0000000110" => data <= "11111111";
            when d"0000000111" => data <= "11111011";
            when d"0000000112" => data <= "10110101";
            when d"0000000113" => data <= "11110111";
            when d"0000000114" => data <= "11111101";
            when d"0000000115" => data <= "11110011";
            when d"0000000116" => data <= "11010111";
            when d"0000000117" => data <= "10000011";
            when d"0000000118" => data <= "10000011";
            when d"0000000119" => data <= "11111011";
            when d"0000000120" => data <= "11000011";
            when d"0000000121" => data <= "10111101";
            when d"0000000122" => data <= "11101111";
            when d"0000000123" => data <= "11111111";
            when d"0000000124" => data <= "11110111";
            when d"0000000125" => data <= "11000001";
            when d"0000000126" => data <= "11110111";
            when d"0000000127" => data <= "11111011";
            when d"0000000128" => data <= "11111111";
            when d"0000000129" => data <= "11101111";
            when d"0000000130" => data <= "11111111";
            when d"0000000131" => data <= "11011011";
            when d"0000000132" => data <= "11000001";
            when d"0000000133" => data <= "11101111";
            when d"0000000134" => data <= "11010101";
            when d"0000000135" => data <= "11111111";
            when d"0000000136" => data <= "11110111";
            when d"0000000137" => data <= "11101111";
            when d"0000000138" => data <= "11000001";
            when d"0000000139" => data <= "11000001";
            when d"0000000140" => data <= "11111111";
            when d"0000000141" => data <= "11000001";
            when d"0000000142" => data <= "11111111";
            when d"0000000143" => data <= "11110111";
            when d"0000000144" => data <= "10101101";
            when d"0000000145" => data <= "11110111";
            when d"0000000146" => data <= "11000011";
            when d"0000000147" => data <= "11111101";
            when d"0000000148" => data <= "10110111";
            when d"0000000149" => data <= "11111101";
            when d"0000000150" => data <= "10111101";
            when d"0000000151" => data <= "11110111";
            when d"0000000152" => data <= "10111101";
            when d"0000000153" => data <= "11000001";
            when d"0000000154" => data <= "11111111";
            when d"0000000155" => data <= "11111111";
            when d"0000000156" => data <= "11101111";
            when d"0000000157" => data <= "11111111";
            when d"0000000158" => data <= "11111011";
            when d"0000000159" => data <= "11110111";
            when d"0000000160" => data <= "11111111";
            when d"0000000161" => data <= "11111111";
            when d"0000000162" => data <= "11111111";
            when d"0000000163" => data <= "10000001";
            when d"0000000164" => data <= "11110101";
            when d"0000000165" => data <= "11011001";
            when d"0000000166" => data <= "10111011";
            when d"0000000167" => data <= "11111111";
            when d"0000000168" => data <= "11110111";
            when d"0000000169" => data <= "11101111";
            when d"0000000170" => data <= "11110111";
            when d"0000000171" => data <= "11110111";
            when d"0000000172" => data <= "11110111";
            when d"0000000173" => data <= "11111111";
            when d"0000000174" => data <= "11100111";
            when d"0000000175" => data <= "11101111";
            when d"0000000176" => data <= "10011101";
            when d"0000000177" => data <= "11110111";
            when d"0000000178" => data <= "10111111";
            when d"0000000179" => data <= "10111101";
            when d"0000000180" => data <= "10000001";
            when d"0000000181" => data <= "10111101";
            when d"0000000182" => data <= "10111101";
            when d"0000000183" => data <= "11101111";
            when d"0000000184" => data <= "10111101";
            when d"0000000185" => data <= "11111101";
            when d"0000000186" => data <= "11111111";
            when d"0000000187" => data <= "11101111";
            when d"0000000188" => data <= "11110111";
            when d"0000000189" => data <= "11000001";
            when d"0000000190" => data <= "11110111";
            when d"0000000191" => data <= "11111111";
            when d"0000000192" => data <= "11111111";
            when d"0000000193" => data <= "11101111";
            when d"0000000194" => data <= "11111111";
            when d"0000000195" => data <= "11011011";
            when d"0000000196" => data <= "11000001";
            when d"0000000197" => data <= "10111001";
            when d"0000000198" => data <= "11000101";
            when d"0000000199" => data <= "11111111";
            when d"0000000200" => data <= "11111011";
            when d"0000000201" => data <= "11011111";
            when d"0000000202" => data <= "11101011";
            when d"0000000203" => data <= "11110111";
            when d"0000000204" => data <= "11110111";
            when d"0000000205" => data <= "11111111";
            when d"0000000206" => data <= "11100111";
            when d"0000000207" => data <= "11011111";
            when d"0000000208" => data <= "11000011";
            when d"0000000209" => data <= "11000001";
            when d"0000000210" => data <= "10000001";
            when d"0000000211" => data <= "11000011";
            when d"0000000212" => data <= "11110111";
            when d"0000000213" => data <= "11000011";
            when d"0000000214" => data <= "11000011";
            when d"0000000215" => data <= "11101111";
            when d"0000000216" => data <= "11000011";
            when d"0000000217" => data <= "11000011";
            when d"0000000218" => data <= "11101111";
            when d"0000000219" => data <= "11101111";
            when d"0000000220" => data <= "11111011";
            when d"0000000221" => data <= "11111111";
            when d"0000000222" => data <= "11101111";
            when d"0000000223" => data <= "11110111";
            when d"0000000224" => data <= "11111111";
            when d"0000000225" => data <= "11111111";
            when d"0000000226" => data <= "11111111";
            when d"0000000227" => data <= "11111111";
            when d"0000000228" => data <= "11110111";
            when d"0000000229" => data <= "11111111";
            when d"0000000230" => data <= "11111111";
            when d"0000000231" => data <= "11111111";
            when d"0000000232" => data <= "11111111";
            when d"0000000233" => data <= "11111111";
            when d"0000000234" => data <= "11111111";
            when d"0000000235" => data <= "11111111";
            when d"0000000236" => data <= "11101111";
            when d"0000000237" => data <= "11111111";
            when d"0000000238" => data <= "11111111";
            when d"0000000239" => data <= "11111111";
            when d"0000000240" => data <= "11111111";
            when d"0000000241" => data <= "11111111";
            when d"0000000242" => data <= "11111111";
            when d"0000000243" => data <= "11111111";
            when d"0000000244" => data <= "11111111";
            when d"0000000245" => data <= "11111111";
            when d"0000000246" => data <= "11111111";
            when d"0000000247" => data <= "11111111";
            when d"0000000248" => data <= "11111111";
            when d"0000000249" => data <= "11111111";
            when d"0000000250" => data <= "11111111";
            when d"0000000251" => data <= "11011111";
            when d"0000000252" => data <= "11111111";
            when d"0000000253" => data <= "11111111";
            when d"0000000254" => data <= "11111111";
            when d"0000000255" => data <= "11111111";
            when d"0000000256" => data <= "11111111";
            when d"0000000257" => data <= "11111111";
            when d"0000000258" => data <= "11111111";
            when d"0000000259" => data <= "11111111";
            when d"0000000260" => data <= "11111111";
            when d"0000000261" => data <= "11111111";
            when d"0000000262" => data <= "11111111";
            when d"0000000263" => data <= "11111111";
            when d"0000000264" => data <= "11111111";
            when d"0000000265" => data <= "11111111";
            when d"0000000266" => data <= "11111111";
            when d"0000000267" => data <= "11111111";
            when d"0000000268" => data <= "11111111";
            when d"0000000269" => data <= "11111111";
            when d"0000000270" => data <= "11111111";
            when d"0000000271" => data <= "11111111";
            when d"0000000272" => data <= "11111111";
            when d"0000000273" => data <= "11111111";
            when d"0000000274" => data <= "11111111";
            when d"0000000275" => data <= "11111111";
            when d"0000000276" => data <= "11111111";
            when d"0000000277" => data <= "11111111";
            when d"0000000278" => data <= "11111111";
            when d"0000000279" => data <= "11111111";
            when d"0000000280" => data <= "11111111";
            when d"0000000281" => data <= "11111111";
            when d"0000000282" => data <= "11111111";
            when d"0000000283" => data <= "11111111";
            when d"0000000284" => data <= "11111111";
            when d"0000000285" => data <= "11111111";
            when d"0000000286" => data <= "11111111";
            when d"0000000287" => data <= "11111111";
            when d"0000000288" => data <= "11000011";
            when d"0000000289" => data <= "11000011";
            when d"0000000290" => data <= "10000011";
            when d"0000000291" => data <= "11000011";
            when d"0000000292" => data <= "10000111";
            when d"0000000293" => data <= "10000001";
            when d"0000000294" => data <= "10000001";
            when d"0000000295" => data <= "11000011";
            when d"0000000296" => data <= "10111101";
            when d"0000000297" => data <= "11000001";
            when d"0000000298" => data <= "11111101";
            when d"0000000299" => data <= "10111011";
            when d"0000000300" => data <= "10111111";
            when d"0000000301" => data <= "10111101";
            when d"0000000302" => data <= "10111101";
            when d"0000000303" => data <= "11000011";
            when d"0000000304" => data <= "10000011";
            when d"0000000305" => data <= "11000011";
            when d"0000000306" => data <= "10000011";
            when d"0000000307" => data <= "11000011";
            when d"0000000308" => data <= "00000001";
            when d"0000000309" => data <= "10111101";
            when d"0000000310" => data <= "10111101";
            when d"0000000311" => data <= "10111101";
            when d"0000000312" => data <= "10111101";
            when d"0000000313" => data <= "01111101";
            when d"0000000314" => data <= "10000001";
            when d"0000000315" => data <= "11110001";
            when d"0000000316" => data <= "11111111";
            when d"0000000317" => data <= "10001111";
            when d"0000000318" => data <= "11101111";
            when d"0000000319" => data <= "11111111";
            when d"0000000320" => data <= "10110101";
            when d"0000000321" => data <= "10111101";
            when d"0000000322" => data <= "10111101";
            when d"0000000323" => data <= "10111101";
            when d"0000000324" => data <= "10111011";
            when d"0000000325" => data <= "10111111";
            when d"0000000326" => data <= "10111111";
            when d"0000000327" => data <= "10111101";
            when d"0000000328" => data <= "10111101";
            when d"0000000329" => data <= "11110111";
            when d"0000000330" => data <= "11111101";
            when d"0000000331" => data <= "10110111";
            when d"0000000332" => data <= "10111111";
            when d"0000000333" => data <= "10011001";
            when d"0000000334" => data <= "10011101";
            when d"0000000335" => data <= "10111101";
            when d"0000000336" => data <= "10111101";
            when d"0000000337" => data <= "10111101";
            when d"0000000338" => data <= "10111101";
            when d"0000000339" => data <= "10111111";
            when d"0000000340" => data <= "11101111";
            when d"0000000341" => data <= "10111101";
            when d"0000000342" => data <= "10111101";
            when d"0000000343" => data <= "10111101";
            when d"0000000344" => data <= "11011011";
            when d"0000000345" => data <= "10111011";
            when d"0000000346" => data <= "11111011";
            when d"0000000347" => data <= "11110111";
            when d"0000000348" => data <= "10111111";
            when d"0000000349" => data <= "11101111";
            when d"0000000350" => data <= "11000111";
            when d"0000000351" => data <= "11111111";
            when d"0000000352" => data <= "10101001";
            when d"0000000353" => data <= "10111101";
            when d"0000000354" => data <= "10000011";
            when d"0000000355" => data <= "10111111";
            when d"0000000356" => data <= "10111101";
            when d"0000000357" => data <= "10000011";
            when d"0000000358" => data <= "10000011";
            when d"0000000359" => data <= "10111111";
            when d"0000000360" => data <= "10000001";
            when d"0000000361" => data <= "11110111";
            when d"0000000362" => data <= "11111101";
            when d"0000000363" => data <= "10001111";
            when d"0000000364" => data <= "10111111";
            when d"0000000365" => data <= "10100101";
            when d"0000000366" => data <= "10101101";
            when d"0000000367" => data <= "10111101";
            when d"0000000368" => data <= "10111101";
            when d"0000000369" => data <= "10111101";
            when d"0000000370" => data <= "10111101";
            when d"0000000371" => data <= "11000011";
            when d"0000000372" => data <= "11101111";
            when d"0000000373" => data <= "10111101";
            when d"0000000374" => data <= "10111101";
            when d"0000000375" => data <= "10111101";
            when d"0000000376" => data <= "11100111";
            when d"0000000377" => data <= "11010111";
            when d"0000000378" => data <= "11110111";
            when d"0000000379" => data <= "11110111";
            when d"0000000380" => data <= "11011111";
            when d"0000000381" => data <= "11101111";
            when d"0000000382" => data <= "10101011";
            when d"0000000383" => data <= "11111111";
            when d"0000000384" => data <= "10100001";
            when d"0000000385" => data <= "10000001";
            when d"0000000386" => data <= "10111101";
            when d"0000000387" => data <= "10111111";
            when d"0000000388" => data <= "10111101";
            when d"0000000389" => data <= "10111111";
            when d"0000000390" => data <= "10111111";
            when d"0000000391" => data <= "10110001";
            when d"0000000392" => data <= "10111101";
            when d"0000000393" => data <= "11110111";
            when d"0000000394" => data <= "10111101";
            when d"0000000395" => data <= "10110111";
            when d"0000000396" => data <= "10111111";
            when d"0000000397" => data <= "10111101";
            when d"0000000398" => data <= "10110101";
            when d"0000000399" => data <= "10111101";
            when d"0000000400" => data <= "10000011";
            when d"0000000401" => data <= "10101101";
            when d"0000000402" => data <= "10000011";
            when d"0000000403" => data <= "11111101";
            when d"0000000404" => data <= "11101111";
            when d"0000000405" => data <= "10111101";
            when d"0000000406" => data <= "10111101";
            when d"0000000407" => data <= "10111101";
            when d"0000000408" => data <= "11100111";
            when d"0000000409" => data <= "11101111";
            when d"0000000410" => data <= "11101111";
            when d"0000000411" => data <= "11110111";
            when d"0000000412" => data <= "11101111";
            when d"0000000413" => data <= "11101111";
            when d"0000000414" => data <= "11101111";
            when d"0000000415" => data <= "11111111";
            when d"0000000416" => data <= "10111111";
            when d"0000000417" => data <= "10111101";
            when d"0000000418" => data <= "10111101";
            when d"0000000419" => data <= "10111101";
            when d"0000000420" => data <= "10111011";
            when d"0000000421" => data <= "10111111";
            when d"0000000422" => data <= "10111111";
            when d"0000000423" => data <= "10111101";
            when d"0000000424" => data <= "10111101";
            when d"0000000425" => data <= "11110111";
            when d"0000000426" => data <= "10111101";
            when d"0000000427" => data <= "10111011";
            when d"0000000428" => data <= "10111111";
            when d"0000000429" => data <= "10111101";
            when d"0000000430" => data <= "10111001";
            when d"0000000431" => data <= "10111101";
            when d"0000000432" => data <= "10111111";
            when d"0000000433" => data <= "10110101";
            when d"0000000434" => data <= "10111011";
            when d"0000000435" => data <= "10111101";
            when d"0000000436" => data <= "11101111";
            when d"0000000437" => data <= "10111101";
            when d"0000000438" => data <= "11011011";
            when d"0000000439" => data <= "10100101";
            when d"0000000440" => data <= "11011011";
            when d"0000000441" => data <= "11101111";
            when d"0000000442" => data <= "11011111";
            when d"0000000443" => data <= "11110111";
            when d"0000000444" => data <= "11110111";
            when d"0000000445" => data <= "11101111";
            when d"0000000446" => data <= "11101111";
            when d"0000000447" => data <= "11111111";
            when d"0000000448" => data <= "11000011";
            when d"0000000449" => data <= "10111101";
            when d"0000000450" => data <= "10000011";
            when d"0000000451" => data <= "11000011";
            when d"0000000452" => data <= "10000111";
            when d"0000000453" => data <= "10000001";
            when d"0000000454" => data <= "10111111";
            when d"0000000455" => data <= "11000011";
            when d"0000000456" => data <= "10111101";
            when d"0000000457" => data <= "11000001";
            when d"0000000458" => data <= "11000011";
            when d"0000000459" => data <= "10111101";
            when d"0000000460" => data <= "10000001";
            when d"0000000461" => data <= "10111101";
            when d"0000000462" => data <= "10111101";
            when d"0000000463" => data <= "11000011";
            when d"0000000464" => data <= "10111111";
            when d"0000000465" => data <= "11000011";
            when d"0000000466" => data <= "10111101";
            when d"0000000467" => data <= "11000011";
            when d"0000000468" => data <= "11101111";
            when d"0000000469" => data <= "11000011";
            when d"0000000470" => data <= "11100111";
            when d"0000000471" => data <= "11011011";
            when d"0000000472" => data <= "10111101";
            when d"0000000473" => data <= "11101111";
            when d"0000000474" => data <= "10000001";
            when d"0000000475" => data <= "11110001";
            when d"0000000476" => data <= "11111111";
            when d"0000000477" => data <= "10001111";
            when d"0000000478" => data <= "11101111";
            when d"0000000479" => data <= "00000000";
            when d"0000000480" => data <= "11111111";
            when d"0000000481" => data <= "11111111";
            when d"0000000482" => data <= "11111111";
            when d"0000000483" => data <= "11111111";
            when d"0000000484" => data <= "11111111";
            when d"0000000485" => data <= "11111111";
            when d"0000000486" => data <= "11111111";
            when d"0000000487" => data <= "11111111";
            when d"0000000488" => data <= "11111111";
            when d"0000000489" => data <= "11111111";
            when d"0000000490" => data <= "11111111";
            when d"0000000491" => data <= "11111111";
            when d"0000000492" => data <= "11111111";
            when d"0000000493" => data <= "11111111";
            when d"0000000494" => data <= "11111111";
            when d"0000000495" => data <= "11111111";
            when d"0000000496" => data <= "11111111";
            when d"0000000497" => data <= "11111111";
            when d"0000000498" => data <= "11111111";
            when d"0000000499" => data <= "11111111";
            when d"0000000500" => data <= "11111111";
            when d"0000000501" => data <= "11111111";
            when d"0000000502" => data <= "11111111";
            when d"0000000503" => data <= "11111111";
            when d"0000000504" => data <= "11111111";
            when d"0000000505" => data <= "11111111";
            when d"0000000506" => data <= "11111111";
            when d"0000000507" => data <= "11111111";
            when d"0000000508" => data <= "11111111";
            when d"0000000509" => data <= "11111111";
            when d"0000000510" => data <= "11111111";
            when d"0000000511" => data <= "11111111";
            when d"0000000512" => data <= "11111111";
            when d"0000000513" => data <= "11111111";
            when d"0000000514" => data <= "11111111";
            when d"0000000515" => data <= "11111111";
            when d"0000000516" => data <= "11111111";
            when d"0000000517" => data <= "11111111";
            when d"0000000518" => data <= "11111111";
            when d"0000000519" => data <= "11111111";
            when d"0000000520" => data <= "11111111";
            when d"0000000521" => data <= "11111111";
            when d"0000000522" => data <= "11111111";
            when d"0000000523" => data <= "11111111";
            when d"0000000524" => data <= "11111111";
            when d"0000000525" => data <= "11111111";
            when d"0000000526" => data <= "11111111";
            when d"0000000527" => data <= "11111111";
            when d"0000000528" => data <= "11111111";
            when d"0000000529" => data <= "11111111";
            when d"0000000530" => data <= "11111111";
            when d"0000000531" => data <= "11111111";
            when d"0000000532" => data <= "11111111";
            when d"0000000533" => data <= "11111111";
            when d"0000000534" => data <= "11111111";
            when d"0000000535" => data <= "11111111";
            when d"0000000536" => data <= "11111111";
            when d"0000000537" => data <= "11111111";
            when d"0000000538" => data <= "11111111";
            when d"0000000539" => data <= "11111111";
            when d"0000000540" => data <= "11111111";
            when d"0000000541" => data <= "11111111";
            when d"0000000542" => data <= "11111111";
            when d"0000000543" => data <= "11000011";
            when d"0000000544" => data <= "11100011";
            when d"0000000545" => data <= "11111111";
            when d"0000000546" => data <= "11011111";
            when d"0000000547" => data <= "11111111";
            when d"0000000548" => data <= "11111011";
            when d"0000000549" => data <= "11111111";
            when d"0000000550" => data <= "11110011";
            when d"0000000551" => data <= "11111111";
            when d"0000000552" => data <= "10111111";
            when d"0000000553" => data <= "11101111";
            when d"0000000554" => data <= "11111011";
            when d"0000000555" => data <= "11011111";
            when d"0000000556" => data <= "11101111";
            when d"0000000557" => data <= "11111111";
            when d"0000000558" => data <= "11111111";
            when d"0000000559" => data <= "11111111";
            when d"0000000560" => data <= "11111111";
            when d"0000000561" => data <= "11111111";
            when d"0000000562" => data <= "11111111";
            when d"0000000563" => data <= "11111111";
            when d"0000000564" => data <= "11101111";
            when d"0000000565" => data <= "11111111";
            when d"0000000566" => data <= "11111111";
            when d"0000000567" => data <= "11111111";
            when d"0000000568" => data <= "11111111";
            when d"0000000569" => data <= "11111111";
            when d"0000000570" => data <= "11111111";
            when d"0000000571" => data <= "11110001";
            when d"0000000572" => data <= "11110111";
            when d"0000000573" => data <= "10001111";
            when d"0000000574" => data <= "11101011";
            when d"0000000575" => data <= "10111101";
            when d"0000000576" => data <= "11011101";
            when d"0000000577" => data <= "11000111";
            when d"0000000578" => data <= "11011111";
            when d"0000000579" => data <= "11100011";
            when d"0000000580" => data <= "11111011";
            when d"0000000581" => data <= "11000111";
            when d"0000000582" => data <= "11101111";
            when d"0000000583" => data <= "11000011";
            when d"0000000584" => data <= "10111111";
            when d"0000000585" => data <= "11111111";
            when d"0000000586" => data <= "11111111";
            when d"0000000587" => data <= "11010111";
            when d"0000000588" => data <= "11101111";
            when d"0000000589" => data <= "10010111";
            when d"0000000590" => data <= "10000111";
            when d"0000000591" => data <= "11000111";
            when d"0000000592" => data <= "10000111";
            when d"0000000593" => data <= "11000011";
            when d"0000000594" => data <= "11100011";
            when d"0000000595" => data <= "11000111";
            when d"0000000596" => data <= "11000111";
            when d"0000000597" => data <= "10111011";
            when d"0000000598" => data <= "10111011";
            when d"0000000599" => data <= "10111011";
            when d"0000000600" => data <= "10111011";
            when d"0000000601" => data <= "10111011";
            when d"0000000602" => data <= "10000011";
            when d"0000000603" => data <= "11110111";
            when d"0000000604" => data <= "11110111";
            when d"0000000605" => data <= "11101111";
            when d"0000000606" => data <= "11010111";
            when d"0000000607" => data <= "01100110";
            when d"0000000608" => data <= "10000111";
            when d"0000000609" => data <= "11111011";
            when d"0000000610" => data <= "11000011";
            when d"0000000611" => data <= "11011111";
            when d"0000000612" => data <= "11000011";
            when d"0000000613" => data <= "10111011";
            when d"0000000614" => data <= "11100111";
            when d"0000000615" => data <= "10111011";
            when d"0000000616" => data <= "10000111";
            when d"0000000617" => data <= "11001111";
            when d"0000000618" => data <= "11111011";
            when d"0000000619" => data <= "11001111";
            when d"0000000620" => data <= "11101111";
            when d"0000000621" => data <= "10101011";
            when d"0000000622" => data <= "10111011";
            when d"0000000623" => data <= "10111011";
            when d"0000000624" => data <= "10111011";
            when d"0000000625" => data <= "10111011";
            when d"0000000626" => data <= "11011111";
            when d"0000000627" => data <= "10111111";
            when d"0000000628" => data <= "11101111";
            when d"0000000629" => data <= "10111011";
            when d"0000000630" => data <= "10111011";
            when d"0000000631" => data <= "10101011";
            when d"0000000632" => data <= "11010111";
            when d"0000000633" => data <= "10111011";
            when d"0000000634" => data <= "11110111";
            when d"0000000635" => data <= "11001111";
            when d"0000000636" => data <= "11110111";
            when d"0000000637" => data <= "11110011";
            when d"0000000638" => data <= "11111111";
            when d"0000000639" => data <= "01011110";
            when d"0000000640" => data <= "11011111";
            when d"0000000641" => data <= "11000011";
            when d"0000000642" => data <= "11011101";
            when d"0000000643" => data <= "11011111";
            when d"0000000644" => data <= "10111011";
            when d"0000000645" => data <= "10000111";
            when d"0000000646" => data <= "11101111";
            when d"0000000647" => data <= "10111011";
            when d"0000000648" => data <= "10111011";
            when d"0000000649" => data <= "11101111";
            when d"0000000650" => data <= "11111011";
            when d"0000000651" => data <= "11001111";
            when d"0000000652" => data <= "11101111";
            when d"0000000653" => data <= "10101011";
            when d"0000000654" => data <= "10111011";
            when d"0000000655" => data <= "10111011";
            when d"0000000656" => data <= "10111011";
            when d"0000000657" => data <= "10111011";
            when d"0000000658" => data <= "11011111";
            when d"0000000659" => data <= "11000111";
            when d"0000000660" => data <= "11101111";
            when d"0000000661" => data <= "10111011";
            when d"0000000662" => data <= "11010111";
            when d"0000000663" => data <= "10101011";
            when d"0000000664" => data <= "11101111";
            when d"0000000665" => data <= "10111011";
            when d"0000000666" => data <= "11101111";
            when d"0000000667" => data <= "11110111";
            when d"0000000668" => data <= "11110111";
            when d"0000000669" => data <= "11101111";
            when d"0000000670" => data <= "11111111";
            when d"0000000671" => data <= "01011110";
            when d"0000000672" => data <= "11011111";
            when d"0000000673" => data <= "10111011";
            when d"0000000674" => data <= "11011101";
            when d"0000000675" => data <= "11011111";
            when d"0000000676" => data <= "10111011";
            when d"0000000677" => data <= "10111111";
            when d"0000000678" => data <= "11101111";
            when d"0000000679" => data <= "11000011";
            when d"0000000680" => data <= "10111011";
            when d"0000000681" => data <= "11101111";
            when d"0000000682" => data <= "11111011";
            when d"0000000683" => data <= "11010111";
            when d"0000000684" => data <= "11101111";
            when d"0000000685" => data <= "10101011";
            when d"0000000686" => data <= "10111011";
            when d"0000000687" => data <= "10111011";
            when d"0000000688" => data <= "10000111";
            when d"0000000689" => data <= "11000011";
            when d"0000000690" => data <= "11011111";
            when d"0000000691" => data <= "11111011";
            when d"0000000692" => data <= "11101111";
            when d"0000000693" => data <= "10111011";
            when d"0000000694" => data <= "11010111";
            when d"0000000695" => data <= "10101011";
            when d"0000000696" => data <= "11010111";
            when d"0000000697" => data <= "11000011";
            when d"0000000698" => data <= "11011111";
            when d"0000000699" => data <= "11110111";
            when d"0000000700" => data <= "11110111";
            when d"0000000701" => data <= "11101111";
            when d"0000000702" => data <= "11111111";
            when d"0000000703" => data <= "01100110";
            when d"0000000704" => data <= "10000001";
            when d"0000000705" => data <= "11000011";
            when d"0000000706" => data <= "11000011";
            when d"0000000707" => data <= "11100011";
            when d"0000000708" => data <= "11000011";
            when d"0000000709" => data <= "11000011";
            when d"0000000710" => data <= "11101111";
            when d"0000000711" => data <= "11111011";
            when d"0000000712" => data <= "10111011";
            when d"0000000713" => data <= "11000111";
            when d"0000000714" => data <= "11011011";
            when d"0000000715" => data <= "11011011";
            when d"0000000716" => data <= "11110011";
            when d"0000000717" => data <= "10101011";
            when d"0000000718" => data <= "10111011";
            when d"0000000719" => data <= "11000111";
            when d"0000000720" => data <= "10111111";
            when d"0000000721" => data <= "11111011";
            when d"0000000722" => data <= "11011111";
            when d"0000000723" => data <= "10000111";
            when d"0000000724" => data <= "11110011";
            when d"0000000725" => data <= "11000111";
            when d"0000000726" => data <= "11101111";
            when d"0000000727" => data <= "11010111";
            when d"0000000728" => data <= "10111011";
            when d"0000000729" => data <= "11111011";
            when d"0000000730" => data <= "10000011";
            when d"0000000731" => data <= "11110001";
            when d"0000000732" => data <= "11110111";
            when d"0000000733" => data <= "10001111";
            when d"0000000734" => data <= "11111111";
            when d"0000000735" => data <= "10111101";
            when d"0000000736" => data <= "11111111";
            when d"0000000737" => data <= "11111111";
            when d"0000000738" => data <= "11111111";
            when d"0000000739" => data <= "11111111";
            when d"0000000740" => data <= "11111111";
            when d"0000000741" => data <= "11111111";
            when d"0000000742" => data <= "11111111";
            when d"0000000743" => data <= "11000111";
            when d"0000000744" => data <= "11111111";
            when d"0000000745" => data <= "11111111";
            when d"0000000746" => data <= "11100111";
            when d"0000000747" => data <= "11111111";
            when d"0000000748" => data <= "11111111";
            when d"0000000749" => data <= "11111111";
            when d"0000000750" => data <= "11111111";
            when d"0000000751" => data <= "11111111";
            when d"0000000752" => data <= "10111111";
            when d"0000000753" => data <= "11111001";
            when d"0000000754" => data <= "11111111";
            when d"0000000755" => data <= "11111111";
            when d"0000000756" => data <= "11111111";
            when d"0000000757" => data <= "11111111";
            when d"0000000758" => data <= "11111111";
            when d"0000000759" => data <= "11111111";
            when d"0000000760" => data <= "11111111";
            when d"0000000761" => data <= "11000111";
            when d"0000000762" => data <= "11111111";
            when d"0000000763" => data <= "11111111";
            when d"0000000764" => data <= "11111111";
            when d"0000000765" => data <= "11111111";
            when d"0000000766" => data <= "11111111";
            when d"0000000767" => data <= "11000011";
            when d"0000000768" => data <= "10000000";
            when d"0000000769" => data <= "01111000";
            when d"0000000770" => data <= "00000111";
            when d"0000000771" => data <= "11111111";
            when d"0000000772" => data <= "10000000";
            when d"0000000773" => data <= "01111000";
            when d"0000000774" => data <= "00000111";
            when d"0000000775" => data <= "11111111";
            when d"0000000776" => data <= "10000000";
            when d"0000000777" => data <= "01111000";
            when d"0000000778" => data <= "00000111";
            when d"0000000779" => data <= "11111111";
            when d"0000000780" => data <= "10000000";
            when d"0000000781" => data <= "01111000";
            when d"0000000782" => data <= "00000111";
            when d"0000000783" => data <= "11111111";
            when d"0000000784" => data <= "11111111";
            when d"0000000785" => data <= "11111111";
            when d"0000000786" => data <= "11111111";
            when d"0000000787" => data <= "11111111";
            when d"0000000788" => data <= "11111111";
            when d"0000000789" => data <= "11111111";
            when d"0000000790" => data <= "11111111";
            when d"0000000791" => data <= "11111111";
            when d"0000000792" => data <= "11111111";
            when d"0000000793" => data <= "11111111";
            when d"0000000794" => data <= "11111111";
            when d"0000000795" => data <= "11111111";
            when d"0000000796" => data <= "11111111";
            when d"0000000797" => data <= "11111111";
            when d"0000000798" => data <= "11111111";
            when d"0000000799" => data <= "11111111";
            when d"0000000800" => data <= "10000000";
            when d"0000000801" => data <= "01111000";
            when d"0000000802" => data <= "00000111";
            when d"0000000803" => data <= "11111111";
            when d"0000000804" => data <= "10000000";
            when d"0000000805" => data <= "01111000";
            when d"0000000806" => data <= "00000111";
            when d"0000000807" => data <= "11111111";
            when d"0000000808" => data <= "10000000";
            when d"0000000809" => data <= "01111000";
            when d"0000000810" => data <= "00000111";
            when d"0000000811" => data <= "11111111";
            when d"0000000812" => data <= "10000000";
            when d"0000000813" => data <= "01111000";
            when d"0000000814" => data <= "00000111";
            when d"0000000815" => data <= "11111111";
            when d"0000000816" => data <= "11111111";
            when d"0000000817" => data <= "11111111";
            when d"0000000818" => data <= "11111111";
            when d"0000000819" => data <= "11111111";
            when d"0000000820" => data <= "11111111";
            when d"0000000821" => data <= "11111111";
            when d"0000000822" => data <= "11111111";
            when d"0000000823" => data <= "11111111";
            when d"0000000824" => data <= "11111111";
            when d"0000000825" => data <= "11111111";
            when d"0000000826" => data <= "11111111";
            when d"0000000827" => data <= "11111111";
            when d"0000000828" => data <= "11111111";
            when d"0000000829" => data <= "11111111";
            when d"0000000830" => data <= "11111111";
            when d"0000000831" => data <= "11111111";
            when d"0000000832" => data <= "10000000";
            when d"0000000833" => data <= "01111000";
            when d"0000000834" => data <= "00000111";
            when d"0000000835" => data <= "11111111";
            when d"0000000836" => data <= "10000000";
            when d"0000000837" => data <= "01111000";
            when d"0000000838" => data <= "00000111";
            when d"0000000839" => data <= "11111111";
            when d"0000000840" => data <= "10000000";
            when d"0000000841" => data <= "01111000";
            when d"0000000842" => data <= "00000111";
            when d"0000000843" => data <= "11111111";
            when d"0000000844" => data <= "10000000";
            when d"0000000845" => data <= "01111000";
            when d"0000000846" => data <= "00000111";
            when d"0000000847" => data <= "11111111";
            when d"0000000848" => data <= "11111111";
            when d"0000000849" => data <= "11111111";
            when d"0000000850" => data <= "11111111";
            when d"0000000851" => data <= "11111111";
            when d"0000000852" => data <= "11111111";
            when d"0000000853" => data <= "11111111";
            when d"0000000854" => data <= "11111111";
            when d"0000000855" => data <= "11111111";
            when d"0000000856" => data <= "11111111";
            when d"0000000857" => data <= "11111111";
            when d"0000000858" => data <= "11111111";
            when d"0000000859" => data <= "11111111";
            when d"0000000860" => data <= "11111111";
            when d"0000000861" => data <= "11111111";
            when d"0000000862" => data <= "11111111";
            when d"0000000863" => data <= "11111111";
            when d"0000000864" => data <= "10000000";
            when d"0000000865" => data <= "01111000";
            when d"0000000866" => data <= "00000111";
            when d"0000000867" => data <= "11111111";
            when d"0000000868" => data <= "10000000";
            when d"0000000869" => data <= "01111000";
            when d"0000000870" => data <= "00000111";
            when d"0000000871" => data <= "11111111";
            when d"0000000872" => data <= "10000000";
            when d"0000000873" => data <= "01111000";
            when d"0000000874" => data <= "00000111";
            when d"0000000875" => data <= "11111111";
            when d"0000000876" => data <= "10000000";
            when d"0000000877" => data <= "01111000";
            when d"0000000878" => data <= "00000111";
            when d"0000000879" => data <= "11111111";
            when d"0000000880" => data <= "11111111";
            when d"0000000881" => data <= "11111111";
            when d"0000000882" => data <= "11111111";
            when d"0000000883" => data <= "11111111";
            when d"0000000884" => data <= "11111111";
            when d"0000000885" => data <= "11111111";
            when d"0000000886" => data <= "11111111";
            when d"0000000887" => data <= "11111111";
            when d"0000000888" => data <= "11111111";
            when d"0000000889" => data <= "11111111";
            when d"0000000890" => data <= "11111111";
            when d"0000000891" => data <= "11111111";
            when d"0000000892" => data <= "11111111";
            when d"0000000893" => data <= "11111111";
            when d"0000000894" => data <= "11111111";
            when d"0000000895" => data <= "11111111";
            when d"0000000896" => data <= "11111111";
            when d"0000000897" => data <= "11111111";
            when d"0000000898" => data <= "11111111";
            when d"0000000899" => data <= "10000111";
            when d"0000000900" => data <= "10000111";
            when d"0000000901" => data <= "10000111";
            when d"0000000902" => data <= "10000000";
            when d"0000000903" => data <= "01111000";
            when d"0000000904" => data <= "01111000";
            when d"0000000905" => data <= "01111000";
            when d"0000000906" => data <= "01111000";
            when d"0000000907" => data <= "00000000";
            when d"0000000908" => data <= "00000000";
            when d"0000000909" => data <= "00000000";
            when d"0000000910" => data <= "00000111";
            when d"0000000911" => data <= "11111111";
            when d"0000000912" => data <= "11111111";
            when d"0000000913" => data <= "11111111";
            when d"0000000914" => data <= "11111111";
            when d"0000000915" => data <= "11111111";
            when d"0000000916" => data <= "11111111";
            when d"0000000917" => data <= "11111111";
            when d"0000000918" => data <= "11111111";
            when d"0000000919" => data <= "11111111";
            when d"0000000920" => data <= "11111111";
            when d"0000000921" => data <= "11111111";
            when d"0000000922" => data <= "11111111";
            when d"0000000923" => data <= "11111111";
            when d"0000000924" => data <= "11111111";
            when d"0000000925" => data <= "11111111";
            when d"0000000926" => data <= "11111111";
            when d"0000000927" => data <= "11111111";
            when d"0000000928" => data <= "11111111";
            when d"0000000929" => data <= "11111111";
            when d"0000000930" => data <= "11111111";
            when d"0000000931" => data <= "10000111";
            when d"0000000932" => data <= "10000111";
            when d"0000000933" => data <= "10000111";
            when d"0000000934" => data <= "10000000";
            when d"0000000935" => data <= "01111000";
            when d"0000000936" => data <= "01111000";
            when d"0000000937" => data <= "01111000";
            when d"0000000938" => data <= "01111000";
            when d"0000000939" => data <= "00000000";
            when d"0000000940" => data <= "00000000";
            when d"0000000941" => data <= "00000000";
            when d"0000000942" => data <= "00000111";
            when d"0000000943" => data <= "11111111";
            when d"0000000944" => data <= "11111111";
            when d"0000000945" => data <= "11111111";
            when d"0000000946" => data <= "11111111";
            when d"0000000947" => data <= "11111111";
            when d"0000000948" => data <= "11111111";
            when d"0000000949" => data <= "11111111";
            when d"0000000950" => data <= "11111111";
            when d"0000000951" => data <= "11111111";
            when d"0000000952" => data <= "11111111";
            when d"0000000953" => data <= "11111111";
            when d"0000000954" => data <= "11111111";
            when d"0000000955" => data <= "11111111";
            when d"0000000956" => data <= "11111111";
            when d"0000000957" => data <= "11111111";
            when d"0000000958" => data <= "11111111";
            when d"0000000959" => data <= "11111111";
            when d"0000000960" => data <= "11111111";
            when d"0000000961" => data <= "11111111";
            when d"0000000962" => data <= "11111111";
            when d"0000000963" => data <= "10000111";
            when d"0000000964" => data <= "10000111";
            when d"0000000965" => data <= "10000111";
            when d"0000000966" => data <= "10000000";
            when d"0000000967" => data <= "01111000";
            when d"0000000968" => data <= "01111000";
            when d"0000000969" => data <= "01111000";
            when d"0000000970" => data <= "01111000";
            when d"0000000971" => data <= "00000000";
            when d"0000000972" => data <= "00000000";
            when d"0000000973" => data <= "00000000";
            when d"0000000974" => data <= "00000111";
            when d"0000000975" => data <= "11111111";
            when d"0000000976" => data <= "11111111";
            when d"0000000977" => data <= "11111111";
            when d"0000000978" => data <= "11111111";
            when d"0000000979" => data <= "11111111";
            when d"0000000980" => data <= "11111111";
            when d"0000000981" => data <= "11111111";
            when d"0000000982" => data <= "11111111";
            when d"0000000983" => data <= "11111111";
            when d"0000000984" => data <= "11111111";
            when d"0000000985" => data <= "11111111";
            when d"0000000986" => data <= "11111111";
            when d"0000000987" => data <= "11111111";
            when d"0000000988" => data <= "11111111";
            when d"0000000989" => data <= "11111111";
            when d"0000000990" => data <= "11111111";
            when d"0000000991" => data <= "11111111";
            when d"0000000992" => data <= "11111111";
            when d"0000000993" => data <= "11111111";
            when d"0000000994" => data <= "11111111";
            when d"0000000995" => data <= "10000111";
            when d"0000000996" => data <= "10000111";
            when d"0000000997" => data <= "10000111";
            when d"0000000998" => data <= "10000000";
            when d"0000000999" => data <= "01111000";
            when d"0000001000" => data <= "01111000";
            when d"0000001001" => data <= "01111000";
            when d"0000001002" => data <= "01111000";
            when d"0000001003" => data <= "00000000";
            when d"0000001004" => data <= "00000000";
            when d"0000001005" => data <= "00000000";
            when d"0000001006" => data <= "00000111";
            when d"0000001007" => data <= "11111111";
            when d"0000001008" => data <= "11111111";
            when d"0000001009" => data <= "11111111";
            when d"0000001010" => data <= "11111111";
            when d"0000001011" => data <= "11111111";
            when d"0000001012" => data <= "11111111";
            when d"0000001013" => data <= "11111111";
            when d"0000001014" => data <= "11111111";
            when d"0000001015" => data <= "11111111";
            when d"0000001016" => data <= "11111111";
            when d"0000001017" => data <= "11111111";
            when d"0000001018" => data <= "11111111";
            when d"0000001019" => data <= "11111111";
            when d"0000001020" => data <= "11111111";
            when d"0000001021" => data <= "11111111";
            when d"0000001022" => data <= "11111111";
            when d"0000001023" => data <= "11111111";
            when others => data <= (others => '0');
        end case;
    end process;
end rtl;
