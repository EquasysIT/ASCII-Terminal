--------------------------------------------------------------
-- Engineer: A Burgess                                      --
--                                                          --
-- Design Name: Computer System ROM                         --
--                                                          --
-- October 2024                                             --
--------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity rom is
	port (
		clk     : in    std_logic;
		addr    : in    std_logic_vector(13 downto 0);
		data    : out   std_logic_vector(7 downto 0)
	);
end;

architecture rtl of rom is
	type romdata is array(0 to 16383) of std_logic_vector(7 downto 0);
	constant rom : romdata := (
		x"4C",x"16",x"DF",x"FB",x"C6",x"08",x"C6",x"16", -- 0x0000
		x"CB",x"B7",x"C7",x"DD",x"C9",x"F0",x"CD",x"09", -- 0x0008
		x"CA",x"64",x"C8",x"64",x"C7",x"3C",x"C7",x"E7", -- 0x0010
		x"C7",x"DD",x"C6",x"47",x"C7",x"91",x"C7",x"FA", -- 0x0018
		x"C7",x"F9",x"C6",x"0A",x"C8",x"6A",x"D5",x"26", -- 0x0020
		x"FF",x"27",x"FF",x"FF",x"D0",x"61",x"D5",x"F3", -- 0x0028
		x"C8",x"22",x"C7",x"79",x"C5",x"3E",x"C5",x"CE", -- 0x0030
		x"C9",x"22",x"C5",x"77",x"D9",x"0A",x"DA",x"96", -- 0x0038
		x"D9",x"00",x"00",x"CC",x"D0",x"ED",x"D0",x"74", -- 0x0040
		x"DC",x"95",x"DD",x"28",x"D7",x"F0",x"DC",x"D1", -- 0x0048
		x"DD",x"D8",x"DD",x"21",x"DE",x"85",x"DE",x"57", -- 0x0050
		x"D5",x"C5",x"D4",x"B2",x"D1",x"F6",x"D4",x"D4", -- 0x0058
		x"D4",x"35",x"D4",x"49",x"D4",x"75",x"D4",x"80", -- 0x0060
		x"D4",x"79",x"A7",x"D5",x"79",x"90",x"D5",x"7B", -- 0x0068
		x"68",x"D7",x"7B",x"4F",x"D8",x"7F",x"7D",x"DC", -- 0x0070
		x"50",x"58",x"CD",x"46",x"55",x"CD",x"7D",x"B6", -- 0x0078
		x"DC",x"5A",x"B2",x"CC",x"64",x"85",x"CD",x"45", -- 0x0080
		x"4E",x"C4",x"46",x"4F",x"D2",x"4E",x"45",x"58", -- 0x0088
		x"D4",x"44",x"41",x"54",x"C1",x"49",x"4E",x"50", -- 0x0090
		x"55",x"D4",x"44",x"49",x"CD",x"52",x"45",x"41", -- 0x0098
		x"C4",x"4C",x"45",x"D4",x"47",x"4F",x"54",x"CF", -- 0x00A0
		x"52",x"55",x"CE",x"49",x"C6",x"52",x"45",x"53", -- 0x00A8
		x"54",x"4F",x"52",x"C5",x"47",x"4F",x"53",x"55", -- 0x00B0
		x"C2",x"52",x"45",x"54",x"55",x"52",x"CE",x"52", -- 0x00B8
		x"45",x"CD",x"53",x"54",x"4F",x"D0",x"4F",x"CE", -- 0x00C0
		x"57",x"41",x"49",x"D4",x"4C",x"4F",x"41",x"C4", -- 0x00C8
		x"53",x"41",x"56",x"C5",x"44",x"45",x"C6",x"50", -- 0x00D0
		x"4F",x"4B",x"C5",x"50",x"52",x"49",x"4E",x"D4", -- 0x00D8
		x"43",x"4F",x"4E",x"D4",x"4C",x"49",x"53",x"D4", -- 0x00E0
		x"43",x"4C",x"45",x"41",x"D2",x"47",x"45",x"D4", -- 0x00E8
		x"4E",x"45",x"D7",x"54",x"41",x"42",x"A8",x"54", -- 0x00F0
		x"CF",x"46",x"CE",x"53",x"50",x"43",x"A8",x"54", -- 0x00F8
		x"48",x"45",x"CE",x"4E",x"4F",x"D4",x"53",x"54", -- 0x0100
		x"45",x"D0",x"AB",x"AD",x"AA",x"AF",x"DE",x"41", -- 0x0108
		x"4E",x"C4",x"4F",x"D2",x"BE",x"BD",x"BC",x"53", -- 0x0110
		x"47",x"CE",x"49",x"4E",x"D4",x"41",x"42",x"D3", -- 0x0118
		x"55",x"53",x"D2",x"46",x"52",x"C5",x"50",x"4F", -- 0x0120
		x"D3",x"53",x"51",x"D2",x"52",x"4E",x"C4",x"4C", -- 0x0128
		x"4F",x"C7",x"45",x"58",x"D0",x"43",x"4F",x"D3", -- 0x0130
		x"53",x"49",x"CE",x"54",x"41",x"CE",x"41",x"54", -- 0x0138
		x"CE",x"50",x"45",x"45",x"CB",x"4C",x"45",x"CE", -- 0x0140
		x"53",x"54",x"52",x"A4",x"56",x"41",x"CC",x"41", -- 0x0148
		x"53",x"C3",x"43",x"48",x"52",x"A4",x"4C",x"45", -- 0x0150
		x"46",x"54",x"A4",x"52",x"49",x"47",x"48",x"54", -- 0x0158
		x"A4",x"4D",x"49",x"44",x"A4",x"47",x"CF",x"00", -- 0x0160
		x"4E",x"45",x"58",x"54",x"20",x"57",x"49",x"54", -- 0x0168
		x"48",x"4F",x"55",x"54",x"20",x"46",x"4F",x"D2", -- 0x0170
		x"53",x"59",x"4E",x"54",x"41",x"D8",x"52",x"45", -- 0x0178
		x"54",x"55",x"52",x"4E",x"20",x"57",x"49",x"54", -- 0x0180
		x"48",x"4F",x"55",x"54",x"20",x"47",x"4F",x"53", -- 0x0188
		x"55",x"C2",x"4F",x"55",x"54",x"20",x"4F",x"46", -- 0x0190
		x"20",x"44",x"41",x"54",x"C1",x"49",x"4C",x"4C", -- 0x0198
		x"45",x"47",x"41",x"4C",x"20",x"51",x"55",x"41", -- 0x01A0
		x"4E",x"54",x"49",x"54",x"D9",x"4F",x"56",x"45", -- 0x01A8
		x"52",x"46",x"4C",x"4F",x"D7",x"4F",x"55",x"54", -- 0x01B0
		x"20",x"4F",x"46",x"20",x"4D",x"45",x"4D",x"4F", -- 0x01B8
		x"52",x"D9",x"55",x"4E",x"44",x"45",x"46",x"27", -- 0x01C0
		x"44",x"20",x"53",x"54",x"41",x"54",x"45",x"4D", -- 0x01C8
		x"45",x"4E",x"D4",x"42",x"41",x"44",x"20",x"53", -- 0x01D0
		x"55",x"42",x"53",x"43",x"52",x"49",x"50",x"D4", -- 0x01D8
		x"52",x"45",x"44",x"49",x"4D",x"27",x"44",x"20", -- 0x01E0
		x"41",x"52",x"52",x"41",x"D9",x"44",x"49",x"56", -- 0x01E8
		x"49",x"53",x"49",x"4F",x"4E",x"20",x"42",x"59", -- 0x01F0
		x"20",x"5A",x"45",x"52",x"CF",x"49",x"4C",x"4C", -- 0x01F8
		x"45",x"47",x"41",x"4C",x"20",x"44",x"49",x"52", -- 0x0200
		x"45",x"43",x"D4",x"54",x"59",x"50",x"45",x"20", -- 0x0208
		x"4D",x"49",x"53",x"4D",x"41",x"54",x"43",x"C8", -- 0x0210
		x"53",x"54",x"52",x"49",x"4E",x"47",x"20",x"54", -- 0x0218
		x"4F",x"4F",x"20",x"4C",x"4F",x"4E",x"C7",x"46", -- 0x0220
		x"4F",x"52",x"4D",x"55",x"4C",x"41",x"20",x"54", -- 0x0228
		x"4F",x"4F",x"20",x"43",x"4F",x"4D",x"50",x"4C", -- 0x0230
		x"45",x"D8",x"43",x"41",x"4E",x"27",x"54",x"20", -- 0x0238
		x"43",x"4F",x"4E",x"54",x"49",x"4E",x"55",x"C5", -- 0x0240
		x"55",x"4E",x"44",x"45",x"46",x"27",x"44",x"20", -- 0x0248
		x"46",x"55",x"4E",x"43",x"54",x"49",x"4F",x"CE", -- 0x0250
		x"20",x"45",x"52",x"52",x"4F",x"52",x"00",x"20", -- 0x0258
		x"49",x"4E",x"20",x"00",x"0D",x"0A",x"4F",x"4B", -- 0x0260
		x"0D",x"0A",x"00",x"0D",x"0A",x"42",x"52",x"45", -- 0x0268
		x"41",x"4B",x"00",x"BA",x"E8",x"E8",x"E8",x"E8", -- 0x0270
		x"BD",x"01",x"01",x"C9",x"81",x"D0",x"21",x"A5", -- 0x0278
		x"9F",x"D0",x"0A",x"BD",x"02",x"01",x"85",x"9E", -- 0x0280
		x"BD",x"03",x"01",x"85",x"9F",x"DD",x"03",x"01", -- 0x0288
		x"D0",x"07",x"A5",x"9E",x"DD",x"02",x"01",x"F0", -- 0x0290
		x"07",x"8A",x"18",x"69",x"12",x"AA",x"D0",x"D8", -- 0x0298
		x"60",x"20",x"F1",x"C2",x"85",x"86",x"84",x"87", -- 0x02A0
		x"38",x"A5",x"AF",x"E5",x"B4",x"85",x"77",x"A8", -- 0x02A8
		x"A5",x"B0",x"E5",x"B5",x"AA",x"E8",x"98",x"F0", -- 0x02B0
		x"23",x"A5",x"AF",x"38",x"E5",x"77",x"85",x"AF", -- 0x02B8
		x"B0",x"03",x"C6",x"B0",x"38",x"A5",x"AD",x"E5", -- 0x02C0
		x"77",x"85",x"AD",x"B0",x"08",x"C6",x"AE",x"90", -- 0x02C8
		x"04",x"B1",x"AF",x"91",x"AD",x"88",x"D0",x"F9", -- 0x02D0
		x"B1",x"AF",x"91",x"AD",x"C6",x"B0",x"C6",x"AE", -- 0x02D8
		x"CA",x"D0",x"F2",x"60",x"0A",x"69",x"3E",x"B0", -- 0x02E0
		x"35",x"85",x"77",x"BA",x"E4",x"77",x"90",x"2E", -- 0x02E8
		x"60",x"C4",x"89",x"90",x"28",x"D0",x"04",x"C5", -- 0x02F0
		x"88",x"90",x"22",x"48",x"A2",x"09",x"98",x"48", -- 0x02F8
		x"B5",x"AC",x"CA",x"10",x"FA",x"20",x"6F",x"D2", -- 0x0300
		x"A2",x"F7",x"68",x"95",x"B6",x"E8",x"30",x"FA", -- 0x0308
		x"68",x"A8",x"68",x"C4",x"89",x"90",x"06",x"D0", -- 0x0310
		x"05",x"C5",x"88",x"B0",x"01",x"60",x"A2",x"4D", -- 0x0318
		x"46",x"6A",x"20",x"32",x"C9",x"20",x"98",x"C9", -- 0x0320
		x"BD",x"68",x"C1",x"48",x"29",x"7F",x"20",x"9A", -- 0x0328
		x"C9",x"E8",x"68",x"10",x"F3",x"20",x"58",x"C5", -- 0x0330
		x"A9",x"58",x"A0",x"C2",x"20",x"78",x"C9",x"A4", -- 0x0338
		x"8F",x"C8",x"F0",x"03",x"20",x"00",x"DB",x"46", -- 0x0340
		x"6A",x"A9",x"64",x"A0",x"C2",x"20",x"03",x"00", -- 0x0348
		x"20",x"28",x"C4",x"86",x"CF",x"84",x"D0",x"20", -- 0x0350
		x"C8",x"00",x"AA",x"F0",x"F3",x"A2",x"FF",x"86", -- 0x0358
		x"8F",x"90",x"06",x"20",x"68",x"C4",x"4C",x"A5", -- 0x0360
		x"C6",x"20",x"2B",x"C8",x"20",x"68",x"C4",x"84", -- 0x0368
		x"62",x"20",x"F4",x"C4",x"90",x"44",x"A0",x"01", -- 0x0370
		x"B1",x"B4",x"85",x"78",x"A5",x"82",x"85",x"77", -- 0x0378
		x"A5",x"B5",x"85",x"7A",x"A5",x"B4",x"88",x"F1", -- 0x0380
		x"B4",x"18",x"65",x"82",x"85",x"82",x"85",x"79", -- 0x0388
		x"A5",x"83",x"69",x"FF",x"85",x"83",x"E5",x"B5", -- 0x0390
		x"AA",x"38",x"A5",x"B4",x"E5",x"82",x"A8",x"B0", -- 0x0398
		x"03",x"E8",x"C6",x"7A",x"18",x"65",x"77",x"90", -- 0x03A0
		x"03",x"C6",x"78",x"18",x"B1",x"77",x"91",x"79", -- 0x03A8
		x"C8",x"D0",x"F9",x"E6",x"78",x"E6",x"7A",x"CA", -- 0x03B0
		x"D0",x"F2",x"20",x"3A",x"C5",x"20",x"F5",x"C3", -- 0x03B8
		x"A5",x"10",x"F0",x"8C",x"18",x"A5",x"82",x"85", -- 0x03C0
		x"AF",x"65",x"62",x"85",x"AD",x"A4",x"83",x"84", -- 0x03C8
		x"B0",x"90",x"01",x"C8",x"84",x"AE",x"20",x"A1", -- 0x03D0
		x"C2",x"A5",x"86",x"A4",x"87",x"85",x"82",x"84", -- 0x03D8
		x"83",x"A4",x"62",x"88",x"B9",x"0C",x"00",x"91", -- 0x03E0
		x"B4",x"88",x"10",x"F8",x"20",x"3A",x"C5",x"20", -- 0x03E8
		x"F5",x"C3",x"4C",x"50",x"C3",x"A5",x"80",x"A4", -- 0x03F0
		x"81",x"85",x"77",x"84",x"78",x"18",x"A0",x"01", -- 0x03F8
		x"B1",x"77",x"F0",x"1D",x"A0",x"04",x"C8",x"B1", -- 0x0400
		x"77",x"D0",x"FB",x"C8",x"98",x"65",x"77",x"AA", -- 0x0408
		x"A0",x"00",x"91",x"77",x"A5",x"78",x"69",x"00", -- 0x0410
		x"C8",x"91",x"77",x"86",x"77",x"85",x"78",x"90", -- 0x0418
		x"DD",x"60",x"CA",x"10",x"05",x"20",x"32",x"C9", -- 0x0420
		x"A2",x"00",x"20",x"58",x"C4",x"C9",x"07",x"F0", -- 0x0428
		x"14",x"C9",x"0D",x"F0",x"20",x"C9",x"20",x"90", -- 0x0430
		x"F1",x"C9",x"7D",x"B0",x"ED",x"C9",x"40",x"F0", -- 0x0438
		x"E4",x"C9",x"5F",x"F0",x"DD",x"E0",x"47",x"B0", -- 0x0440
		x"05",x"95",x"10",x"E8",x"D0",x"DC",x"A9",x"07", -- 0x0448
		x"20",x"9A",x"C9",x"D0",x"D5",x"4C",x"2C",x"C9", -- 0x0450
		x"20",x"07",x"FF",x"C9",x"0F",x"D0",x"08",x"48", -- 0x0458
		x"A5",x"6A",x"49",x"FF",x"85",x"6A",x"68",x"60", -- 0x0460
		x"A6",x"CF",x"A0",x"04",x"84",x"66",x"BD",x"00", -- 0x0468
		x"00",x"C9",x"20",x"F0",x"37",x"85",x"61",x"C9", -- 0x0470
		x"22",x"F0",x"56",x"24",x"66",x"70",x"2D",x"C9", -- 0x0478
		x"3F",x"D0",x"04",x"A9",x"96",x"D0",x"25",x"C9", -- 0x0480
		x"30",x"90",x"04",x"C9",x"3C",x"90",x"1D",x"84", -- 0x0488
		x"C6",x"A0",x"00",x"84",x"62",x"88",x"86",x"CF", -- 0x0490
		x"CA",x"C8",x"E8",x"BD",x"00",x"00",x"38",x"F9", -- 0x0498
		x"87",x"C0",x"F0",x"F5",x"C9",x"80",x"D0",x"30", -- 0x04A0
		x"05",x"62",x"A4",x"C6",x"E8",x"C8",x"99",x"0B", -- 0x04A8
		x"00",x"B9",x"0B",x"00",x"F0",x"36",x"38",x"E9", -- 0x04B0
		x"3A",x"F0",x"04",x"C9",x"49",x"D0",x"02",x"85", -- 0x04B8
		x"66",x"38",x"E9",x"54",x"D0",x"A8",x"85",x"61", -- 0x04C0
		x"BD",x"00",x"00",x"F0",x"DF",x"C5",x"61",x"F0", -- 0x04C8
		x"DB",x"C8",x"99",x"0B",x"00",x"E8",x"D0",x"F0", -- 0x04D0
		x"A6",x"CF",x"E6",x"62",x"C8",x"B9",x"86",x"C0", -- 0x04D8
		x"10",x"FA",x"B9",x"87",x"C0",x"D0",x"B4",x"BD", -- 0x04E0
		x"00",x"00",x"10",x"BE",x"99",x"0D",x"00",x"A9", -- 0x04E8
		x"0F",x"85",x"CF",x"60",x"A5",x"80",x"A6",x"81", -- 0x04F0
		x"A0",x"01",x"85",x"B4",x"86",x"B5",x"B1",x"B4", -- 0x04F8
		x"F0",x"1F",x"C8",x"C8",x"A5",x"0F",x"D1",x"B4", -- 0x0500
		x"90",x"18",x"F0",x"03",x"88",x"D0",x"09",x"A5", -- 0x0508
		x"0E",x"88",x"D1",x"B4",x"90",x"0C",x"F0",x"0A", -- 0x0510
		x"88",x"B1",x"B4",x"AA",x"88",x"B1",x"B4",x"B0", -- 0x0518
		x"D7",x"18",x"60",x"D0",x"FD",x"A9",x"00",x"A8", -- 0x0520
		x"91",x"80",x"C8",x"91",x"80",x"A5",x"80",x"18", -- 0x0528
		x"69",x"02",x"85",x"82",x"A5",x"81",x"69",x"00", -- 0x0530
		x"85",x"83",x"20",x"6C",x"C5",x"A9",x"00",x"D0", -- 0x0538
		x"2A",x"A5",x"8C",x"A4",x"8D",x"85",x"88",x"84", -- 0x0540
		x"89",x"A5",x"82",x"A4",x"83",x"85",x"84",x"84", -- 0x0548
		x"85",x"85",x"86",x"84",x"87",x"20",x"DE",x"C6", -- 0x0550
		x"A2",x"6E",x"86",x"6B",x"68",x"A8",x"68",x"A2", -- 0x0558
		x"FA",x"9A",x"48",x"98",x"48",x"A9",x"00",x"85", -- 0x0560
		x"93",x"85",x"67",x"60",x"18",x"A5",x"80",x"69", -- 0x0568
		x"FF",x"85",x"CF",x"A5",x"81",x"69",x"FF",x"85", -- 0x0570
		x"D0",x"60",x"90",x"06",x"F0",x"04",x"C9",x"A4", -- 0x0578
		x"D0",x"E9",x"20",x"2B",x"C8",x"20",x"F4",x"C4", -- 0x0580
		x"20",x"CE",x"00",x"F0",x"0C",x"C9",x"A4",x"D0", -- 0x0588
		x"91",x"20",x"C8",x"00",x"20",x"2B",x"C8",x"D0", -- 0x0590
		x"89",x"68",x"68",x"A5",x"0E",x"05",x"0F",x"D0", -- 0x0598
		x"06",x"A9",x"FF",x"85",x"0E",x"85",x"0F",x"A0", -- 0x05A0
		x"01",x"B1",x"B4",x"F0",x"39",x"20",x"ED",x"C6", -- 0x05A8
		x"20",x"32",x"C9",x"C8",x"B1",x"B4",x"AA",x"C8", -- 0x05B0
		x"B1",x"B4",x"C5",x"0F",x"D0",x"04",x"E4",x"0E", -- 0x05B8
		x"F0",x"02",x"B0",x"22",x"84",x"9E",x"20",x"0B", -- 0x05C0
		x"DB",x"A9",x"20",x"A4",x"9E",x"29",x"7F",x"20", -- 0x05C8
		x"9A",x"C9",x"C8",x"F0",x"11",x"B1",x"B4",x"D0", -- 0x05D0
		x"10",x"A8",x"B1",x"B4",x"AA",x"C8",x"B1",x"B4", -- 0x05D8
		x"86",x"B4",x"85",x"B5",x"D0",x"C1",x"4C",x"47", -- 0x05E0
		x"C3",x"10",x"E4",x"38",x"E9",x"7F",x"AA",x"84", -- 0x05E8
		x"9E",x"A0",x"FF",x"CA",x"F0",x"08",x"C8",x"B9", -- 0x05F0
		x"87",x"C0",x"10",x"FA",x"30",x"F5",x"C8",x"B9", -- 0x05F8
		x"87",x"C0",x"30",x"C7",x"20",x"9A",x"C9",x"D0", -- 0x0600
		x"F5",x"A9",x"80",x"85",x"67",x"20",x"65",x"C8", -- 0x0608
		x"20",x"73",x"C2",x"D0",x"05",x"8A",x"69",x"0F", -- 0x0610
		x"AA",x"9A",x"68",x"68",x"A9",x"09",x"20",x"E4", -- 0x0618
		x"C2",x"20",x"C6",x"C7",x"18",x"98",x"65",x"CF", -- 0x0620
		x"48",x"A5",x"D0",x"69",x"00",x"48",x"A5",x"8F", -- 0x0628
		x"48",x"A5",x"8E",x"48",x"A9",x"9D",x"20",x"DE", -- 0x0630
		x"CC",x"20",x"85",x"CB",x"20",x"82",x"CB",x"A5", -- 0x0638
		x"BB",x"09",x"7F",x"25",x"B7",x"85",x"B7",x"A9", -- 0x0640
		x"52",x"A0",x"C6",x"85",x"77",x"84",x"78",x"4C", -- 0x0648
		x"3B",x"CC",x"A9",x"FA",x"A0",x"D6",x"20",x"E0", -- 0x0650
		x"D8",x"20",x"CE",x"00",x"C9",x"A2",x"D0",x"06", -- 0x0658
		x"20",x"C8",x"00",x"20",x"82",x"CB",x"20",x"69", -- 0x0660
		x"D9",x"20",x"30",x"CC",x"A5",x"9F",x"48",x"A5", -- 0x0668
		x"9E",x"48",x"A9",x"81",x"48",x"20",x"ED",x"C6", -- 0x0670
		x"A5",x"CF",x"A4",x"D0",x"F0",x"06",x"85",x"92", -- 0x0678
		x"84",x"93",x"A0",x"00",x"B1",x"CF",x"D0",x"40", -- 0x0680
		x"A0",x"02",x"B1",x"CF",x"18",x"D0",x"03",x"4C", -- 0x0688
		x"13",x"C7",x"C8",x"B1",x"CF",x"85",x"8E",x"C8", -- 0x0690
		x"B1",x"CF",x"85",x"8F",x"98",x"65",x"CF",x"85", -- 0x0698
		x"CF",x"90",x"02",x"E6",x"D0",x"20",x"C8",x"00", -- 0x06A0
		x"20",x"AE",x"C6",x"4C",x"75",x"C6",x"F0",x"3C", -- 0x06A8
		x"E9",x"80",x"90",x"11",x"C9",x"1C",x"B0",x"17", -- 0x06B0
		x"0A",x"A8",x"B9",x"04",x"C0",x"48",x"B9",x"03", -- 0x06B8
		x"C0",x"48",x"4C",x"C8",x"00",x"4C",x"65",x"C8", -- 0x06C0
		x"C9",x"3A",x"F0",x"D9",x"4C",x"E7",x"CC",x"C9", -- 0x06C8
		x"44",x"D0",x"F9",x"20",x"C8",x"00",x"A9",x"9D", -- 0x06D0
		x"20",x"DE",x"CC",x"4C",x"65",x"C7",x"38",x"A5", -- 0x06D8
		x"80",x"E9",x"01",x"A4",x"81",x"B0",x"01",x"88", -- 0x06E0
		x"85",x"96",x"84",x"97",x"60",x"20",x"07",x"FF", -- 0x06E8
		x"90",x"07",x"C9",x"03",x"D0",x"03",x"4C",x"FA", -- 0x06F0
		x"C6",x"60",x"B0",x"01",x"18",x"D0",x"3D",x"A5", -- 0x06F8
		x"CF",x"A4",x"D0",x"F0",x"0C",x"85",x"92",x"84", -- 0x0700
		x"93",x"A5",x"8E",x"A4",x"8F",x"85",x"90",x"84", -- 0x0708
		x"91",x"68",x"68",x"A9",x"6B",x"A0",x"C2",x"A2", -- 0x0710
		x"00",x"86",x"6A",x"90",x"03",x"4C",x"3C",x"C3", -- 0x0718
		x"4C",x"47",x"C3",x"D0",x"17",x"A2",x"D2",x"A4", -- 0x0720
		x"93",x"D0",x"03",x"4C",x"20",x"C3",x"A5",x"92", -- 0x0728
		x"85",x"CF",x"84",x"D0",x"A5",x"90",x"A4",x"91", -- 0x0730
		x"85",x"8E",x"84",x"8F",x"60",x"D0",x"03",x"4C", -- 0x0738
		x"3A",x"C5",x"20",x"41",x"C5",x"4C",x"5C",x"C7", -- 0x0740
		x"A9",x"03",x"20",x"E4",x"C2",x"A5",x"D0",x"48", -- 0x0748
		x"A5",x"CF",x"48",x"A5",x"8F",x"48",x"A5",x"8E", -- 0x0750
		x"48",x"A9",x"8C",x"48",x"20",x"CE",x"00",x"20", -- 0x0758
		x"65",x"C7",x"4C",x"75",x"C6",x"20",x"2B",x"C8", -- 0x0760
		x"20",x"C9",x"C7",x"A5",x"8F",x"C5",x"0F",x"B0", -- 0x0768
		x"0B",x"98",x"38",x"65",x"CF",x"A6",x"D0",x"90", -- 0x0770
		x"07",x"E8",x"B0",x"04",x"A5",x"80",x"A6",x"81", -- 0x0778
		x"20",x"F8",x"C4",x"90",x"1E",x"A5",x"B4",x"E9", -- 0x0780
		x"01",x"85",x"CF",x"A5",x"B5",x"E9",x"00",x"85", -- 0x0788
		x"D0",x"60",x"D0",x"FD",x"A9",x"FF",x"85",x"9F", -- 0x0790
		x"20",x"73",x"C2",x"9A",x"C9",x"8C",x"F0",x"0B", -- 0x0798
		x"A2",x"16",x"2C",x"A2",x"5A",x"4C",x"20",x"C3", -- 0x07A0
		x"4C",x"E7",x"CC",x"68",x"68",x"85",x"8E",x"68", -- 0x07A8
		x"85",x"8F",x"68",x"85",x"CF",x"68",x"85",x"D0", -- 0x07B0
		x"20",x"C6",x"C7",x"98",x"18",x"65",x"CF",x"85", -- 0x07B8
		x"CF",x"90",x"02",x"E6",x"D0",x"60",x"A2",x"3A", -- 0x07C0
		x"2C",x"A2",x"00",x"86",x"60",x"A0",x"00",x"84", -- 0x07C8
		x"61",x"A5",x"61",x"A6",x"60",x"85",x"60",x"86", -- 0x07D0
		x"61",x"B1",x"CF",x"F0",x"E8",x"C5",x"61",x"F0", -- 0x07D8
		x"E4",x"C8",x"C9",x"22",x"D0",x"F3",x"F0",x"E9", -- 0x07E0
		x"20",x"96",x"CB",x"20",x"CE",x"00",x"C9",x"88", -- 0x07E8
		x"F0",x"05",x"A9",x"A0",x"20",x"DE",x"CC",x"A5", -- 0x07F0
		x"B6",x"D0",x"05",x"20",x"C9",x"C7",x"F0",x"BB", -- 0x07F8
		x"20",x"CE",x"00",x"B0",x"03",x"4C",x"65",x"C7", -- 0x0800
		x"4C",x"AE",x"C6",x"20",x"E7",x"D4",x"48",x"C9", -- 0x0808
		x"8C",x"F0",x"04",x"C9",x"88",x"D0",x"91",x"C6", -- 0x0810
		x"BA",x"D0",x"04",x"68",x"4C",x"B0",x"C6",x"20", -- 0x0818
		x"C8",x"00",x"20",x"2B",x"C8",x"C9",x"2C",x"F0", -- 0x0820
		x"EE",x"68",x"60",x"A2",x"00",x"86",x"0E",x"86", -- 0x0828
		x"0F",x"B0",x"F7",x"E9",x"2F",x"85",x"60",x"A5", -- 0x0830
		x"0F",x"85",x"77",x"C9",x"19",x"B0",x"D4",x"A5", -- 0x0838
		x"0E",x"0A",x"26",x"77",x"0A",x"26",x"77",x"65", -- 0x0840
		x"0E",x"85",x"0E",x"A5",x"77",x"65",x"0F",x"85", -- 0x0848
		x"0F",x"06",x"0E",x"26",x"0F",x"A5",x"0E",x"65", -- 0x0850
		x"60",x"85",x"0E",x"90",x"02",x"E6",x"0F",x"20", -- 0x0858
		x"C8",x"00",x"4C",x"31",x"C8",x"20",x"FB",x"CD", -- 0x0860
		x"85",x"9E",x"84",x"9F",x"A9",x"AB",x"20",x"DE", -- 0x0868
		x"CC",x"A5",x"65",x"48",x"A5",x"64",x"48",x"20", -- 0x0870
		x"96",x"CB",x"68",x"2A",x"20",x"88",x"CB",x"D0", -- 0x0878
		x"18",x"68",x"10",x"12",x"20",x"59",x"D9",x"20", -- 0x0880
		x"0D",x"CF",x"A0",x"00",x"A5",x"B9",x"91",x"9E", -- 0x0888
		x"C8",x"A5",x"BA",x"91",x"9E",x"60",x"4C",x"0E", -- 0x0890
		x"D9",x"68",x"A0",x"02",x"B1",x"B9",x"C5",x"89", -- 0x0898
		x"90",x"17",x"D0",x"07",x"88",x"B1",x"B9",x"C5", -- 0x08A0
		x"88",x"90",x"0E",x"A4",x"BA",x"C4",x"83",x"90", -- 0x08A8
		x"08",x"D0",x"0D",x"A5",x"B9",x"C5",x"82",x"B0", -- 0x08B0
		x"07",x"A5",x"B9",x"A4",x"BA",x"4C",x"D6",x"C8", -- 0x08B8
		x"A0",x"00",x"B1",x"B9",x"20",x"C2",x"D1",x"A5", -- 0x08C0
		x"A5",x"A4",x"A6",x"85",x"C4",x"84",x"C5",x"20", -- 0x08C8
		x"C3",x"D3",x"A9",x"B6",x"A0",x"00",x"85",x"A5", -- 0x08D0
		x"84",x"A6",x"20",x"24",x"D4",x"A0",x"00",x"B1", -- 0x08D8
		x"A5",x"91",x"9E",x"C8",x"B1",x"A5",x"91",x"9E", -- 0x08E0
		x"C8",x"B1",x"A5",x"91",x"9E",x"60",x"20",x"7B", -- 0x08E8
		x"C9",x"20",x"CE",x"00",x"F0",x"3C",x"F0",x"48", -- 0x08F0
		x"C9",x"9C",x"F0",x"5C",x"C9",x"9F",x"18",x"F0", -- 0x08F8
		x"57",x"C9",x"2C",x"F0",x"3C",x"C9",x"3B",x"F0", -- 0x0900
		x"64",x"20",x"96",x"CB",x"24",x"64",x"30",x"DE", -- 0x0908
		x"20",x"1B",x"DB",x"20",x"D4",x"D1",x"A0",x"00", -- 0x0910
		x"B1",x"B9",x"18",x"65",x"0B",x"C5",x"0C",x"90", -- 0x0918
		x"03",x"20",x"32",x"C9",x"20",x"7B",x"C9",x"20", -- 0x0920
		x"95",x"C9",x"D0",x"C5",x"A0",x"00",x"94",x"10", -- 0x0928
		x"A2",x"0F",x"A9",x"0D",x"85",x"0B",x"20",x"9A", -- 0x0930
		x"C9",x"A9",x"0A",x"20",x"9A",x"C9",x"49",x"FF", -- 0x0938
		x"60",x"A5",x"0B",x"C5",x"0D",x"90",x"06",x"20", -- 0x0940
		x"32",x"C9",x"4C",x"6D",x"C9",x"38",x"E9",x"0E", -- 0x0948
		x"B0",x"FC",x"49",x"FF",x"69",x"01",x"D0",x"10", -- 0x0950
		x"08",x"20",x"E4",x"D4",x"C9",x"29",x"D0",x"5C", -- 0x0958
		x"28",x"90",x"06",x"8A",x"E5",x"0B",x"90",x"05", -- 0x0960
		x"AA",x"E8",x"CA",x"D0",x"06",x"20",x"C8",x"00", -- 0x0968
		x"4C",x"F6",x"C8",x"20",x"95",x"C9",x"D0",x"F2", -- 0x0970
		x"20",x"D4",x"D1",x"20",x"EF",x"D3",x"AA",x"A0", -- 0x0978
		x"00",x"E8",x"CA",x"F0",x"BB",x"B1",x"77",x"20", -- 0x0980
		x"9A",x"C9",x"C8",x"C9",x"0D",x"D0",x"F3",x"20", -- 0x0988
		x"3E",x"C9",x"4C",x"82",x"C9",x"A9",x"20",x"2C", -- 0x0990
		x"A9",x"3F",x"24",x"6A",x"30",x"09",x"C9",x"20", -- 0x0998
		x"90",x"02",x"E6",x"0B",x"20",x"FC",x"FE",x"29", -- 0x09A0
		x"FF",x"60",x"A5",x"68",x"F0",x"11",x"30",x"04", -- 0x09A8
		x"A0",x"FF",x"D0",x"04",x"A5",x"94",x"A4",x"95", -- 0x09B0
		x"85",x"8E",x"84",x"8F",x"4C",x"E7",x"CC",x"A9", -- 0x09B8
		x"04",x"A0",x"CB",x"20",x"78",x"C9",x"A5",x"92", -- 0x09C0
		x"A4",x"93",x"85",x"CF",x"84",x"D0",x"60",x"20", -- 0x09C8
		x"F3",x"D0",x"A2",x"11",x"A0",x"00",x"84",x"11", -- 0x09D0
		x"A9",x"40",x"20",x"10",x"CA",x"60",x"46",x"6A", -- 0x09D8
		x"C9",x"22",x"D0",x"0B",x"20",x"9C",x"CC",x"A9", -- 0x09E0
		x"3B",x"20",x"DE",x"CC",x"20",x"7B",x"C9",x"20", -- 0x09E8
		x"F3",x"D0",x"A9",x"2C",x"85",x"0F",x"20",x"01", -- 0x09F0
		x"CA",x"A5",x"10",x"D0",x"12",x"18",x"4C",x"09", -- 0x09F8
		x"C7",x"20",x"98",x"C9",x"20",x"95",x"C9",x"4C", -- 0x0A00
		x"28",x"C4",x"A6",x"96",x"A4",x"97",x"A9",x"98", -- 0x0A08
		x"85",x"68",x"86",x"98",x"84",x"99",x"20",x"FB", -- 0x0A10
		x"CD",x"85",x"9E",x"84",x"9F",x"A5",x"CF",x"A4", -- 0x0A18
		x"D0",x"85",x"0E",x"84",x"0F",x"A6",x"98",x"A4", -- 0x0A20
		x"99",x"86",x"CF",x"84",x"D0",x"20",x"CE",x"00", -- 0x0A28
		x"D0",x"1B",x"24",x"68",x"50",x"0B",x"20",x"07", -- 0x0A30
		x"FF",x"85",x"10",x"A2",x"0F",x"A0",x"00",x"F0", -- 0x0A38
		x"08",x"30",x"71",x"20",x"98",x"C9",x"20",x"01", -- 0x0A40
		x"CA",x"86",x"CF",x"84",x"D0",x"20",x"C8",x"00", -- 0x0A48
		x"24",x"64",x"10",x"31",x"24",x"68",x"50",x"09", -- 0x0A50
		x"E8",x"86",x"CF",x"A9",x"00",x"85",x"60",x"F0", -- 0x0A58
		x"0C",x"85",x"60",x"C9",x"22",x"F0",x"07",x"A9", -- 0x0A60
		x"3A",x"85",x"60",x"A9",x"2C",x"18",x"85",x"61", -- 0x0A68
		x"A5",x"CF",x"A4",x"D0",x"69",x"00",x"90",x"01", -- 0x0A70
		x"C8",x"20",x"DA",x"D1",x"20",x"2C",x"D5",x"20", -- 0x0A78
		x"9A",x"C8",x"4C",x"8D",x"CA",x"20",x"31",x"DA", -- 0x0A80
		x"A5",x"65",x"20",x"82",x"C8",x"20",x"CE",x"00", -- 0x0A88
		x"F0",x"07",x"C9",x"2C",x"F0",x"03",x"4C",x"AA", -- 0x0A90
		x"C9",x"A5",x"CF",x"A4",x"D0",x"85",x"98",x"84", -- 0x0A98
		x"99",x"A5",x"0E",x"A4",x"0F",x"85",x"CF",x"84", -- 0x0AA0
		x"D0",x"20",x"CE",x"00",x"F0",x"2C",x"20",x"DC", -- 0x0AA8
		x"CC",x"4C",x"16",x"CA",x"20",x"C6",x"C7",x"C8", -- 0x0AB0
		x"AA",x"D0",x"12",x"A2",x"2A",x"C8",x"B1",x"CF", -- 0x0AB8
		x"F0",x"69",x"C8",x"B1",x"CF",x"85",x"94",x"C8", -- 0x0AC0
		x"B1",x"CF",x"C8",x"85",x"95",x"B1",x"CF",x"AA", -- 0x0AC8
		x"20",x"BB",x"C7",x"E0",x"83",x"D0",x"DD",x"4C", -- 0x0AD0
		x"4D",x"CA",x"A5",x"98",x"A4",x"99",x"A6",x"68", -- 0x0AD8
		x"10",x"03",x"4C",x"E8",x"C6",x"A0",x"00",x"B1", -- 0x0AE0
		x"98",x"F0",x"07",x"A9",x"F3",x"A0",x"CA",x"4C", -- 0x0AE8
		x"78",x"C9",x"60",x"3F",x"45",x"58",x"54",x"52", -- 0x0AF0
		x"41",x"20",x"49",x"47",x"4E",x"4F",x"52",x"45", -- 0x0AF8
		x"44",x"0D",x"0A",x"00",x"3F",x"52",x"45",x"44", -- 0x0B00
		x"4F",x"20",x"46",x"52",x"4F",x"4D",x"20",x"53", -- 0x0B08
		x"54",x"41",x"52",x"54",x"0D",x"0A",x"00",x"D0", -- 0x0B10
		x"04",x"A0",x"00",x"F0",x"03",x"20",x"FB",x"CD", -- 0x0B18
		x"85",x"9E",x"84",x"9F",x"20",x"73",x"C2",x"F0", -- 0x0B20
		x"04",x"A2",x"00",x"F0",x"66",x"9A",x"8A",x"18", -- 0x0B28
		x"69",x"04",x"48",x"69",x"06",x"85",x"79",x"68", -- 0x0B30
		x"A0",x"01",x"20",x"E0",x"D8",x"BA",x"BD",x"09", -- 0x0B38
		x"01",x"85",x"BB",x"A5",x"9E",x"A4",x"9F",x"20", -- 0x0B40
		x"A5",x"D5",x"20",x"0E",x"D9",x"A0",x"01",x"20", -- 0x0B48
		x"9B",x"D9",x"BA",x"38",x"FD",x"09",x"01",x"F0", -- 0x0B50
		x"17",x"BD",x"0F",x"01",x"85",x"8E",x"BD",x"10", -- 0x0B58
		x"01",x"85",x"8F",x"BD",x"12",x"01",x"85",x"CF", -- 0x0B60
		x"BD",x"11",x"01",x"85",x"D0",x"4C",x"75",x"C6", -- 0x0B68
		x"8A",x"69",x"11",x"AA",x"9A",x"20",x"CE",x"00", -- 0x0B70
		x"C9",x"2C",x"D0",x"F1",x"20",x"C8",x"00",x"20", -- 0x0B78
		x"1D",x"CB",x"20",x"96",x"CB",x"18",x"24",x"38", -- 0x0B80
		x"24",x"64",x"30",x"03",x"B0",x"03",x"60",x"B0", -- 0x0B88
		x"FD",x"A2",x"A3",x"4C",x"20",x"C3",x"A6",x"CF", -- 0x0B90
		x"D0",x"02",x"C6",x"D0",x"C6",x"CF",x"A2",x"00", -- 0x0B98
		x"24",x"48",x"8A",x"48",x"A9",x"01",x"20",x"E4", -- 0x0BA0
		x"C2",x"20",x"7B",x"CC",x"A9",x"00",x"85",x"A2", -- 0x0BA8
		x"20",x"CE",x"00",x"38",x"E9",x"AA",x"90",x"17", -- 0x0BB0
		x"C9",x"03",x"B0",x"13",x"C9",x"01",x"2A",x"49", -- 0x0BB8
		x"01",x"45",x"A2",x"C5",x"A2",x"90",x"61",x"85", -- 0x0BC0
		x"A2",x"20",x"C8",x"00",x"4C",x"B3",x"CB",x"A6", -- 0x0BC8
		x"A2",x"D0",x"2C",x"B0",x"7B",x"69",x"07",x"90", -- 0x0BD0
		x"77",x"65",x"64",x"D0",x"03",x"4C",x"86",x"D3", -- 0x0BD8
		x"69",x"FF",x"85",x"77",x"0A",x"65",x"77",x"A8", -- 0x0BE0
		x"68",x"D9",x"69",x"C0",x"B0",x"67",x"20",x"85", -- 0x0BE8
		x"CB",x"48",x"20",x"18",x"CC",x"68",x"A4",x"A0", -- 0x0BF0
		x"10",x"17",x"AA",x"F0",x"56",x"D0",x"5F",x"46", -- 0x0BF8
		x"64",x"8A",x"2A",x"A6",x"CF",x"D0",x"02",x"C6", -- 0x0C00
		x"D0",x"C6",x"CF",x"A0",x"1B",x"85",x"A2",x"D0", -- 0x0C08
		x"D7",x"D9",x"69",x"C0",x"B0",x"48",x"90",x"D9", -- 0x0C10
		x"B9",x"6B",x"C0",x"48",x"B9",x"6A",x"C0",x"48", -- 0x0C18
		x"20",x"2B",x"CC",x"A5",x"A2",x"4C",x"A1",x"CB", -- 0x0C20
		x"4C",x"E7",x"CC",x"A5",x"BB",x"BE",x"69",x"C0", -- 0x0C28
		x"A8",x"68",x"85",x"77",x"E6",x"77",x"68",x"85", -- 0x0C30
		x"78",x"98",x"48",x"20",x"59",x"D9",x"A5",x"BA", -- 0x0C38
		x"48",x"A5",x"B9",x"48",x"A5",x"B8",x"48",x"A5", -- 0x0C40
		x"B7",x"48",x"A5",x"B6",x"48",x"6C",x"77",x"00", -- 0x0C48
		x"A0",x"FF",x"68",x"F0",x"23",x"C9",x"64",x"F0", -- 0x0C50
		x"03",x"20",x"85",x"CB",x"84",x"A0",x"68",x"4A", -- 0x0C58
		x"85",x"69",x"68",x"85",x"BE",x"68",x"85",x"BF", -- 0x0C60
		x"68",x"85",x"C0",x"68",x"85",x"C1",x"68",x"85", -- 0x0C68
		x"C2",x"68",x"85",x"C3",x"45",x"BB",x"85",x"C4", -- 0x0C70
		x"A5",x"B6",x"60",x"A9",x"00",x"85",x"64",x"20", -- 0x0C78
		x"C8",x"00",x"B0",x"03",x"4C",x"31",x"DA",x"20", -- 0x0C80
		x"85",x"CE",x"B0",x"67",x"C9",x"2E",x"F0",x"F4", -- 0x0C88
		x"C9",x"A4",x"F0",x"58",x"C9",x"A3",x"F0",x"E7", -- 0x0C90
		x"C9",x"22",x"D0",x"0F",x"A5",x"CF",x"A4",x"D0", -- 0x0C98
		x"69",x"00",x"90",x"01",x"C8",x"20",x"D4",x"D1", -- 0x0CA0
		x"4C",x"2C",x"D5",x"C9",x"A1",x"D0",x"13",x"A0", -- 0x0CA8
		x"18",x"D0",x"3B",x"20",x"0D",x"CF",x"A5",x"BA", -- 0x0CB0
		x"49",x"FF",x"A8",x"A5",x"B9",x"49",x"FF",x"4C", -- 0x0CB8
		x"E0",x"D0",x"C9",x"9E",x"D0",x"03",x"4C",x"41", -- 0x0CC0
		x"D1",x"C9",x"AD",x"90",x"03",x"4C",x"17",x"CD", -- 0x0CC8
		x"20",x"D9",x"CC",x"20",x"96",x"CB",x"A9",x"29", -- 0x0CD0
		x"2C",x"A9",x"28",x"2C",x"A9",x"2C",x"A0",x"00", -- 0x0CD8
		x"D1",x"CF",x"D0",x"03",x"4C",x"C8",x"00",x"A2", -- 0x0CE0
		x"10",x"4C",x"20",x"C3",x"A0",x"15",x"68",x"68", -- 0x0CE8
		x"4C",x"F2",x"CB",x"20",x"FB",x"CD",x"85",x"B9", -- 0x0CF0
		x"84",x"BA",x"A6",x"64",x"F0",x"05",x"A2",x"00", -- 0x0CF8
		x"86",x"C5",x"60",x"A6",x"65",x"10",x"0D",x"A0", -- 0x0D00
		x"00",x"B1",x"B9",x"AA",x"C8",x"B1",x"B9",x"A8", -- 0x0D08
		x"8A",x"4C",x"E0",x"D0",x"4C",x"E0",x"D8",x"0A", -- 0x0D10
		x"48",x"AA",x"20",x"C8",x"00",x"E0",x"81",x"90", -- 0x0D18
		x"20",x"20",x"D9",x"CC",x"20",x"96",x"CB",x"20", -- 0x0D20
		x"DC",x"CC",x"20",x"87",x"CB",x"68",x"AA",x"A5", -- 0x0D28
		x"BA",x"48",x"A5",x"B9",x"48",x"8A",x"48",x"20", -- 0x0D30
		x"E7",x"D4",x"68",x"A8",x"8A",x"48",x"4C",x"46", -- 0x0D38
		x"CD",x"20",x"D0",x"CC",x"68",x"A8",x"B9",x"E1", -- 0x0D40
		x"BF",x"85",x"AA",x"B9",x"E2",x"BF",x"85",x"AB", -- 0x0D48
		x"20",x"A9",x"00",x"4C",x"85",x"CB",x"A0",x"FF", -- 0x0D50
		x"2C",x"A0",x"00",x"84",x"62",x"20",x"0D",x"CF", -- 0x0D58
		x"A5",x"B9",x"45",x"62",x"85",x"60",x"A5",x"BA", -- 0x0D60
		x"45",x"62",x"85",x"61",x"20",x"3A",x"D9",x"20", -- 0x0D68
		x"0D",x"CF",x"A5",x"BA",x"45",x"62",x"25",x"61", -- 0x0D70
		x"45",x"62",x"A8",x"A5",x"B9",x"45",x"62",x"25", -- 0x0D78
		x"60",x"45",x"62",x"4C",x"E0",x"D0",x"20",x"88", -- 0x0D80
		x"CB",x"B0",x"13",x"A5",x"C3",x"09",x"7F",x"25", -- 0x0D88
		x"BF",x"85",x"BF",x"A9",x"BE",x"A0",x"00",x"20", -- 0x0D90
		x"99",x"D9",x"AA",x"4C",x"D1",x"CD",x"A9",x"00", -- 0x0D98
		x"85",x"64",x"C6",x"A2",x"20",x"EF",x"D3",x"85", -- 0x0DA0
		x"B6",x"86",x"B7",x"84",x"B8",x"A5",x"C1",x"A4", -- 0x0DA8
		x"C2",x"20",x"F3",x"D3",x"86",x"C1",x"84",x"C2", -- 0x0DB0
		x"AA",x"38",x"E5",x"B6",x"F0",x"08",x"A9",x"01", -- 0x0DB8
		x"90",x"04",x"A6",x"B6",x"A9",x"FF",x"85",x"BB", -- 0x0DC0
		x"A0",x"FF",x"E8",x"C8",x"CA",x"D0",x"07",x"A6", -- 0x0DC8
		x"BB",x"30",x"0F",x"18",x"90",x"0C",x"B1",x"C1", -- 0x0DD0
		x"D1",x"B7",x"F0",x"EF",x"A2",x"FF",x"B0",x"02", -- 0x0DD8
		x"A2",x"01",x"E8",x"8A",x"2A",x"25",x"69",x"F0", -- 0x0DE0
		x"02",x"A9",x"FF",x"4C",x"7A",x"D9",x"20",x"DC", -- 0x0DE8
		x"CC",x"AA",x"20",x"00",x"CE",x"20",x"CE",x"00", -- 0x0DF0
		x"D0",x"F4",x"60",x"A2",x"00",x"20",x"CE",x"00", -- 0x0DF8
		x"86",x"63",x"85",x"9A",x"20",x"CE",x"00",x"20", -- 0x0E00
		x"85",x"CE",x"B0",x"03",x"4C",x"E7",x"CC",x"A2", -- 0x0E08
		x"00",x"86",x"64",x"86",x"65",x"20",x"C8",x"00", -- 0x0E10
		x"90",x"05",x"20",x"85",x"CE",x"90",x"0B",x"AA", -- 0x0E18
		x"20",x"C8",x"00",x"90",x"FB",x"20",x"85",x"CE", -- 0x0E20
		x"B0",x"F6",x"C9",x"24",x"D0",x"06",x"A9",x"FF", -- 0x0E28
		x"85",x"64",x"D0",x"10",x"C9",x"25",x"D0",x"13", -- 0x0E30
		x"A5",x"67",x"D0",x"D0",x"A9",x"80",x"85",x"65", -- 0x0E38
		x"05",x"9A",x"85",x"9A",x"8A",x"09",x"80",x"AA", -- 0x0E40
		x"20",x"C8",x"00",x"86",x"9B",x"38",x"05",x"67", -- 0x0E48
		x"E9",x"28",x"D0",x"03",x"4C",x"1F",x"CF",x"A9", -- 0x0E50
		x"00",x"85",x"67",x"A5",x"82",x"A6",x"83",x"A0", -- 0x0E58
		x"00",x"86",x"B5",x"85",x"B4",x"E4",x"85",x"D0", -- 0x0E60
		x"04",x"C5",x"84",x"F0",x"22",x"A5",x"9A",x"D1", -- 0x0E68
		x"B4",x"D0",x"08",x"A5",x"9B",x"C8",x"D1",x"B4", -- 0x0E70
		x"F0",x"62",x"88",x"18",x"A5",x"B4",x"69",x"07", -- 0x0E78
		x"90",x"E1",x"E8",x"D0",x"DC",x"C9",x"41",x"90", -- 0x0E80
		x"05",x"E9",x"5B",x"38",x"E9",x"A5",x"60",x"68", -- 0x0E88
		x"48",x"C9",x"F5",x"D0",x"05",x"A9",x"4D",x"A0", -- 0x0E90
		x"DC",x"60",x"A5",x"84",x"A4",x"85",x"85",x"B4", -- 0x0E98
		x"84",x"B5",x"A5",x"86",x"A4",x"87",x"85",x"AF", -- 0x0EA0
		x"84",x"B0",x"18",x"69",x"07",x"90",x"01",x"C8", -- 0x0EA8
		x"85",x"AD",x"84",x"AE",x"20",x"A1",x"C2",x"A5", -- 0x0EB0
		x"AD",x"A4",x"AE",x"C8",x"85",x"84",x"84",x"85", -- 0x0EB8
		x"A0",x"00",x"A5",x"9A",x"91",x"B4",x"C8",x"A5", -- 0x0EC0
		x"9B",x"91",x"B4",x"A9",x"00",x"C8",x"91",x"B4", -- 0x0EC8
		x"C8",x"91",x"B4",x"C8",x"91",x"B4",x"C8",x"91", -- 0x0ED0
		x"B4",x"C8",x"91",x"B4",x"A5",x"B4",x"18",x"69", -- 0x0ED8
		x"02",x"A4",x"B5",x"90",x"01",x"C8",x"85",x"9C", -- 0x0EE0
		x"84",x"9D",x"60",x"A5",x"62",x"0A",x"69",x"05", -- 0x0EE8
		x"65",x"B4",x"A4",x"B5",x"90",x"01",x"C8",x"85", -- 0x0EF0
		x"AD",x"84",x"AE",x"60",x"90",x"80",x"00",x"00", -- 0x0EF8
		x"20",x"C8",x"00",x"20",x"96",x"CB",x"20",x"85", -- 0x0F00
		x"CB",x"A5",x"BB",x"30",x"0D",x"A5",x"B6",x"C9", -- 0x0F08
		x"90",x"90",x"09",x"A9",x"FC",x"A0",x"CE",x"20", -- 0x0F10
		x"99",x"D9",x"D0",x"7A",x"4C",x"D9",x"D9",x"A5", -- 0x0F18
		x"63",x"05",x"65",x"48",x"A5",x"64",x"48",x"A0", -- 0x0F20
		x"00",x"98",x"48",x"A5",x"9B",x"48",x"A5",x"9A", -- 0x0F28
		x"48",x"20",x"00",x"CF",x"68",x"85",x"9A",x"68", -- 0x0F30
		x"85",x"9B",x"68",x"A8",x"BA",x"BD",x"02",x"01", -- 0x0F38
		x"48",x"BD",x"01",x"01",x"48",x"A5",x"B9",x"9D", -- 0x0F40
		x"02",x"01",x"A5",x"BA",x"9D",x"01",x"01",x"C8", -- 0x0F48
		x"20",x"CE",x"00",x"C9",x"2C",x"F0",x"D2",x"84", -- 0x0F50
		x"62",x"20",x"D6",x"CC",x"68",x"85",x"64",x"68", -- 0x0F58
		x"85",x"65",x"29",x"7F",x"85",x"63",x"A6",x"84", -- 0x0F60
		x"A5",x"85",x"86",x"B4",x"85",x"B5",x"C5",x"87", -- 0x0F68
		x"D0",x"04",x"E4",x"86",x"F0",x"39",x"A0",x"00", -- 0x0F70
		x"B1",x"B4",x"C8",x"C5",x"9A",x"D0",x"06",x"A5", -- 0x0F78
		x"9B",x"D1",x"B4",x"F0",x"16",x"C8",x"B1",x"B4", -- 0x0F80
		x"18",x"65",x"B4",x"AA",x"C8",x"B1",x"B4",x"65", -- 0x0F88
		x"B5",x"90",x"D7",x"A2",x"6B",x"2C",x"A2",x"35", -- 0x0F90
		x"4C",x"20",x"C3",x"A2",x"78",x"A5",x"63",x"D0", -- 0x0F98
		x"F7",x"20",x"EB",x"CE",x"A5",x"62",x"A0",x"04", -- 0x0FA0
		x"D1",x"B4",x"D0",x"E7",x"4C",x"39",x"D0",x"20", -- 0x0FA8
		x"EB",x"CE",x"20",x"F1",x"C2",x"A9",x"00",x"A8", -- 0x0FB0
		x"85",x"C7",x"A2",x"05",x"A5",x"9A",x"91",x"B4", -- 0x0FB8
		x"10",x"01",x"CA",x"C8",x"A5",x"9B",x"91",x"B4", -- 0x0FC0
		x"10",x"02",x"CA",x"CA",x"86",x"C6",x"A5",x"62", -- 0x0FC8
		x"C8",x"C8",x"C8",x"91",x"B4",x"A2",x"0B",x"A9", -- 0x0FD0
		x"00",x"24",x"63",x"50",x"08",x"68",x"18",x"69", -- 0x0FD8
		x"01",x"AA",x"68",x"69",x"00",x"C8",x"91",x"B4", -- 0x0FE0
		x"C8",x"8A",x"91",x"B4",x"20",x"9B",x"D0",x"86", -- 0x0FE8
		x"C6",x"85",x"C7",x"A4",x"77",x"C6",x"62",x"D0", -- 0x0FF0
		x"DC",x"65",x"AE",x"B0",x"5D",x"85",x"AE",x"A8", -- 0x0FF8
		x"8A",x"65",x"AD",x"90",x"03",x"C8",x"F0",x"52", -- 0x1000
		x"20",x"F1",x"C2",x"85",x"86",x"84",x"87",x"A9", -- 0x1008
		x"00",x"E6",x"C7",x"A4",x"C6",x"F0",x"05",x"88", -- 0x1010
		x"91",x"AD",x"D0",x"FB",x"C6",x"AE",x"C6",x"C7", -- 0x1018
		x"D0",x"F5",x"E6",x"AE",x"38",x"A5",x"86",x"E5", -- 0x1020
		x"B4",x"A0",x"02",x"91",x"B4",x"A5",x"87",x"C8", -- 0x1028
		x"E5",x"B5",x"91",x"B4",x"A5",x"63",x"D0",x"62", -- 0x1030
		x"C8",x"B1",x"B4",x"85",x"62",x"A9",x"00",x"85", -- 0x1038
		x"C6",x"85",x"C7",x"C8",x"68",x"AA",x"85",x"B9", -- 0x1040
		x"68",x"85",x"BA",x"D1",x"B4",x"90",x"0E",x"D0", -- 0x1048
		x"06",x"C8",x"8A",x"D1",x"B4",x"90",x"07",x"4C", -- 0x1050
		x"93",x"CF",x"4C",x"1E",x"C3",x"C8",x"A5",x"C7", -- 0x1058
		x"05",x"C6",x"18",x"F0",x"0A",x"20",x"9B",x"D0", -- 0x1060
		x"8A",x"65",x"B9",x"AA",x"98",x"A4",x"77",x"65", -- 0x1068
		x"BA",x"86",x"C6",x"C6",x"62",x"D0",x"CA",x"85", -- 0x1070
		x"C7",x"A2",x"05",x"A5",x"9A",x"10",x"01",x"CA", -- 0x1078
		x"A5",x"9B",x"10",x"02",x"CA",x"CA",x"86",x"7D", -- 0x1080
		x"A9",x"00",x"20",x"A4",x"D0",x"8A",x"65",x"AD", -- 0x1088
		x"85",x"9C",x"98",x"65",x"AE",x"85",x"9D",x"A8", -- 0x1090
		x"A5",x"9C",x"60",x"84",x"77",x"B1",x"B4",x"85", -- 0x1098
		x"7D",x"88",x"B1",x"B4",x"85",x"7E",x"A9",x"10", -- 0x10A0
		x"85",x"B2",x"A2",x"00",x"A0",x"00",x"8A",x"0A", -- 0x10A8
		x"AA",x"98",x"2A",x"A8",x"B0",x"A4",x"06",x"C6", -- 0x10B0
		x"26",x"C7",x"90",x"0B",x"18",x"8A",x"65",x"7D", -- 0x10B8
		x"AA",x"98",x"65",x"7E",x"A8",x"B0",x"93",x"C6", -- 0x10C0
		x"B2",x"D0",x"E3",x"60",x"A5",x"64",x"F0",x"03", -- 0x10C8
		x"20",x"EF",x"D3",x"20",x"6F",x"D2",x"38",x"A5", -- 0x10D0
		x"88",x"E5",x"86",x"A8",x"A5",x"89",x"E5",x"87", -- 0x10D8
		x"A2",x"00",x"86",x"64",x"85",x"B7",x"84",x"B8", -- 0x10E0
		x"A2",x"90",x"4C",x"82",x"D9",x"A4",x"0B",x"A9", -- 0x10E8
		x"00",x"F0",x"ED",x"A6",x"8F",x"E8",x"D0",x"A2", -- 0x10F0
		x"A2",x"95",x"2C",x"A2",x"E0",x"4C",x"20",x"C3", -- 0x10F8
		x"20",x"2E",x"D1",x"20",x"F3",x"D0",x"20",x"D9", -- 0x1100
		x"CC",x"A9",x"80",x"85",x"67",x"20",x"FB",x"CD", -- 0x1108
		x"20",x"85",x"CB",x"20",x"D6",x"CC",x"A9",x"AB", -- 0x1110
		x"20",x"DE",x"CC",x"48",x"A5",x"9D",x"48",x"A5", -- 0x1118
		x"9C",x"48",x"A5",x"D0",x"48",x"A5",x"CF",x"48", -- 0x1120
		x"20",x"B8",x"C7",x"4C",x"9C",x"D1",x"A9",x"9E", -- 0x1128
		x"20",x"DE",x"CC",x"09",x"80",x"85",x"67",x"20", -- 0x1130
		x"02",x"CE",x"85",x"A3",x"84",x"A4",x"4C",x"85", -- 0x1138
		x"CB",x"20",x"2E",x"D1",x"A5",x"A4",x"48",x"A5", -- 0x1140
		x"A3",x"48",x"20",x"D0",x"CC",x"20",x"85",x"CB", -- 0x1148
		x"68",x"85",x"A3",x"68",x"85",x"A4",x"A0",x"02", -- 0x1150
		x"B1",x"A3",x"85",x"9C",x"AA",x"C8",x"B1",x"A3", -- 0x1158
		x"F0",x"99",x"85",x"9D",x"C8",x"B1",x"9C",x"48", -- 0x1160
		x"88",x"10",x"FA",x"A4",x"9D",x"20",x"12",x"D9", -- 0x1168
		x"A5",x"D0",x"48",x"A5",x"CF",x"48",x"B1",x"A3", -- 0x1170
		x"85",x"CF",x"C8",x"B1",x"A3",x"85",x"D0",x"A5", -- 0x1178
		x"9D",x"48",x"A5",x"9C",x"48",x"20",x"82",x"CB", -- 0x1180
		x"68",x"85",x"A3",x"68",x"85",x"A4",x"20",x"CE", -- 0x1188
		x"00",x"F0",x"03",x"4C",x"E7",x"CC",x"68",x"85", -- 0x1190
		x"CF",x"68",x"85",x"D0",x"A0",x"00",x"68",x"91", -- 0x1198
		x"A3",x"68",x"C8",x"91",x"A3",x"68",x"C8",x"91", -- 0x11A0
		x"A3",x"68",x"C8",x"91",x"A3",x"68",x"C8",x"91", -- 0x11A8
		x"A3",x"60",x"20",x"85",x"CB",x"A0",x"00",x"20", -- 0x11B0
		x"1D",x"DB",x"68",x"68",x"A9",x"FF",x"A0",x"00", -- 0x11B8
		x"F0",x"12",x"A6",x"B9",x"A4",x"BA",x"86",x"A5", -- 0x11C0
		x"84",x"A6",x"20",x"3D",x"D2",x"86",x"B7",x"84", -- 0x11C8
		x"B8",x"85",x"B6",x"60",x"A2",x"22",x"86",x"60", -- 0x11D0
		x"86",x"61",x"85",x"C4",x"84",x"C5",x"85",x"B7", -- 0x11D8
		x"84",x"B8",x"A0",x"FF",x"C8",x"B1",x"C4",x"F0", -- 0x11E0
		x"0C",x"C5",x"60",x"F0",x"04",x"C5",x"61",x"D0", -- 0x11E8
		x"F3",x"C9",x"22",x"F0",x"01",x"18",x"84",x"B6", -- 0x11F0
		x"98",x"65",x"C4",x"85",x"C6",x"A6",x"C5",x"90", -- 0x11F8
		x"01",x"E8",x"86",x"C7",x"A5",x"C5",x"D0",x"0B", -- 0x1200
		x"98",x"20",x"C2",x"D1",x"A6",x"C4",x"A4",x"C5", -- 0x1208
		x"20",x"D1",x"D3",x"A6",x"6B",x"E0",x"77",x"D0", -- 0x1210
		x"05",x"A2",x"BF",x"4C",x"20",x"C3",x"A5",x"B6", -- 0x1218
		x"95",x"00",x"A5",x"B7",x"95",x"01",x"A5",x"B8", -- 0x1220
		x"95",x"02",x"A0",x"00",x"86",x"B9",x"84",x"BA", -- 0x1228
		x"84",x"C5",x"88",x"84",x"64",x"86",x"6C",x"E8", -- 0x1230
		x"E8",x"E8",x"86",x"6B",x"60",x"46",x"66",x"48", -- 0x1238
		x"49",x"FF",x"38",x"65",x"88",x"A4",x"89",x"B0", -- 0x1240
		x"01",x"88",x"C4",x"87",x"90",x"11",x"D0",x"04", -- 0x1248
		x"C5",x"86",x"90",x"0B",x"85",x"88",x"84",x"89", -- 0x1250
		x"85",x"8A",x"84",x"8B",x"AA",x"68",x"60",x"A2", -- 0x1258
		x"4D",x"A5",x"66",x"30",x"B6",x"20",x"6F",x"D2", -- 0x1260
		x"A9",x"80",x"85",x"66",x"68",x"D0",x"D0",x"A6", -- 0x1268
		x"8C",x"A5",x"8D",x"86",x"88",x"85",x"89",x"A0", -- 0x1270
		x"00",x"84",x"A4",x"84",x"A3",x"A5",x"86",x"A6", -- 0x1278
		x"87",x"85",x"B4",x"86",x"B5",x"A9",x"6E",x"A2", -- 0x1280
		x"00",x"85",x"77",x"86",x"78",x"C5",x"6B",x"F0", -- 0x1288
		x"05",x"20",x"10",x"D3",x"F0",x"F7",x"A9",x"07", -- 0x1290
		x"85",x"A8",x"A5",x"82",x"A6",x"83",x"85",x"77", -- 0x1298
		x"86",x"78",x"E4",x"85",x"D0",x"04",x"C5",x"84", -- 0x12A0
		x"F0",x"05",x"20",x"06",x"D3",x"F0",x"F3",x"85", -- 0x12A8
		x"AD",x"86",x"AE",x"A9",x"03",x"85",x"A8",x"A5", -- 0x12B0
		x"AD",x"A6",x"AE",x"E4",x"87",x"D0",x"07",x"C5", -- 0x12B8
		x"86",x"D0",x"03",x"4C",x"4F",x"D3",x"85",x"77", -- 0x12C0
		x"86",x"78",x"A0",x"00",x"B1",x"77",x"AA",x"C8", -- 0x12C8
		x"B1",x"77",x"08",x"C8",x"B1",x"77",x"65",x"AD", -- 0x12D0
		x"85",x"AD",x"C8",x"B1",x"77",x"65",x"AE",x"85", -- 0x12D8
		x"AE",x"28",x"10",x"D3",x"8A",x"30",x"D0",x"C8", -- 0x12E0
		x"B1",x"77",x"A0",x"00",x"0A",x"69",x"05",x"65", -- 0x12E8
		x"77",x"85",x"77",x"90",x"02",x"E6",x"78",x"A6", -- 0x12F0
		x"78",x"E4",x"AE",x"D0",x"04",x"C5",x"AD",x"F0", -- 0x12F8
		x"BA",x"20",x"10",x"D3",x"F0",x"F3",x"B1",x"77", -- 0x1300
		x"30",x"35",x"C8",x"B1",x"77",x"10",x"30",x"C8", -- 0x1308
		x"B1",x"77",x"F0",x"2B",x"C8",x"B1",x"77",x"AA", -- 0x1310
		x"C8",x"B1",x"77",x"C5",x"89",x"90",x"06",x"D0", -- 0x1318
		x"1E",x"E4",x"88",x"B0",x"1A",x"C5",x"B5",x"90", -- 0x1320
		x"16",x"D0",x"04",x"E4",x"B4",x"90",x"10",x"86", -- 0x1328
		x"B4",x"85",x"B5",x"A5",x"77",x"A6",x"78",x"85", -- 0x1330
		x"A3",x"86",x"A4",x"A5",x"A8",x"85",x"AA",x"A5", -- 0x1338
		x"A8",x"18",x"65",x"77",x"85",x"77",x"90",x"02", -- 0x1340
		x"E6",x"78",x"A6",x"78",x"A0",x"00",x"60",x"A5", -- 0x1348
		x"A4",x"05",x"A3",x"F0",x"F5",x"A5",x"AA",x"29", -- 0x1350
		x"04",x"4A",x"A8",x"85",x"AA",x"B1",x"A3",x"65", -- 0x1358
		x"B4",x"85",x"AF",x"A5",x"B5",x"69",x"00",x"85", -- 0x1360
		x"B0",x"A5",x"88",x"A6",x"89",x"85",x"AD",x"86", -- 0x1368
		x"AE",x"20",x"A8",x"C2",x"A4",x"AA",x"C8",x"A5", -- 0x1370
		x"AD",x"91",x"A3",x"AA",x"E6",x"AE",x"A5",x"AE", -- 0x1378
		x"C8",x"91",x"A3",x"4C",x"73",x"D2",x"A5",x"BA", -- 0x1380
		x"48",x"A5",x"B9",x"48",x"20",x"7B",x"CC",x"20", -- 0x1388
		x"87",x"CB",x"68",x"85",x"C4",x"68",x"85",x"C5", -- 0x1390
		x"A0",x"00",x"B1",x"C4",x"18",x"71",x"B9",x"90", -- 0x1398
		x"05",x"A2",x"B0",x"4C",x"20",x"C3",x"20",x"C2", -- 0x13A0
		x"D1",x"20",x"C3",x"D3",x"A5",x"A5",x"A4",x"A6", -- 0x13A8
		x"20",x"F3",x"D3",x"20",x"D5",x"D3",x"A5",x"C4", -- 0x13B0
		x"A4",x"C5",x"20",x"F3",x"D3",x"20",x"13",x"D2", -- 0x13B8
		x"4C",x"B0",x"CB",x"A0",x"00",x"B1",x"C4",x"48", -- 0x13C0
		x"C8",x"B1",x"C4",x"AA",x"C8",x"B1",x"C4",x"A8", -- 0x13C8
		x"68",x"86",x"77",x"84",x"78",x"A8",x"F0",x"0A", -- 0x13D0
		x"48",x"88",x"B1",x"77",x"91",x"8A",x"98",x"D0", -- 0x13D8
		x"F8",x"68",x"18",x"65",x"8A",x"85",x"8A",x"90", -- 0x13E0
		x"02",x"E6",x"8B",x"60",x"20",x"87",x"CB",x"A5", -- 0x13E8
		x"B9",x"A4",x"BA",x"85",x"77",x"84",x"78",x"20", -- 0x13F0
		x"24",x"D4",x"08",x"A0",x"00",x"B1",x"77",x"48", -- 0x13F8
		x"C8",x"B1",x"77",x"AA",x"C8",x"B1",x"77",x"A8", -- 0x1400
		x"68",x"28",x"D0",x"13",x"C4",x"89",x"D0",x"0F", -- 0x1408
		x"E4",x"88",x"D0",x"0B",x"48",x"18",x"65",x"88", -- 0x1410
		x"85",x"88",x"90",x"02",x"E6",x"89",x"68",x"86", -- 0x1418
		x"77",x"84",x"78",x"60",x"C4",x"6D",x"D0",x"0C", -- 0x1420
		x"C5",x"6C",x"D0",x"08",x"85",x"6B",x"E9",x"03", -- 0x1428
		x"85",x"6C",x"A0",x"00",x"60",x"20",x"EA",x"D4", -- 0x1430
		x"8A",x"48",x"A9",x"01",x"20",x"CA",x"D1",x"68", -- 0x1438
		x"A0",x"00",x"91",x"B7",x"68",x"68",x"4C",x"13", -- 0x1440
		x"D2",x"20",x"AA",x"D4",x"D1",x"A5",x"98",x"90", -- 0x1448
		x"04",x"B1",x"A5",x"AA",x"98",x"48",x"8A",x"48", -- 0x1450
		x"20",x"CA",x"D1",x"A5",x"A5",x"A4",x"A6",x"20", -- 0x1458
		x"F3",x"D3",x"68",x"A8",x"68",x"18",x"65",x"77", -- 0x1460
		x"85",x"77",x"90",x"02",x"E6",x"78",x"98",x"20", -- 0x1468
		x"D5",x"D3",x"4C",x"13",x"D2",x"20",x"AA",x"D4", -- 0x1470
		x"18",x"F1",x"A5",x"49",x"FF",x"4C",x"4F",x"D4", -- 0x1478
		x"A9",x"FF",x"85",x"BA",x"20",x"CE",x"00",x"C9", -- 0x1480
		x"29",x"F0",x"06",x"20",x"DC",x"CC",x"20",x"E7", -- 0x1488
		x"D4",x"20",x"AA",x"D4",x"F0",x"4B",x"CA",x"8A", -- 0x1490
		x"48",x"18",x"A2",x"00",x"F1",x"A5",x"B0",x"B6", -- 0x1498
		x"49",x"FF",x"C5",x"BA",x"90",x"B1",x"A5",x"BA", -- 0x14A0
		x"B0",x"AD",x"20",x"D6",x"CC",x"68",x"A8",x"68", -- 0x14A8
		x"85",x"AA",x"68",x"68",x"68",x"AA",x"68",x"85", -- 0x14B0
		x"A5",x"68",x"85",x"A6",x"A5",x"AA",x"48",x"98", -- 0x14B8
		x"48",x"A0",x"00",x"8A",x"60",x"20",x"CB",x"D4", -- 0x14C0
		x"4C",x"EF",x"D0",x"20",x"EC",x"D3",x"A2",x"00", -- 0x14C8
		x"86",x"64",x"A8",x"60",x"20",x"CB",x"D4",x"F0", -- 0x14D0
		x"08",x"A0",x"00",x"B1",x"77",x"A8",x"4C",x"EF", -- 0x14D8
		x"D0",x"4C",x"96",x"CF",x"20",x"C8",x"00",x"20", -- 0x14E0
		x"82",x"CB",x"20",x"06",x"CF",x"A6",x"B9",x"D0", -- 0x14E8
		x"F0",x"A6",x"BA",x"4C",x"CE",x"00",x"20",x"CB", -- 0x14F0
		x"D4",x"D0",x"03",x"4C",x"35",x"D6",x"A6",x"CF", -- 0x14F8
		x"A4",x"D0",x"86",x"C6",x"84",x"C7",x"A6",x"77", -- 0x1500
		x"86",x"CF",x"18",x"65",x"77",x"85",x"79",x"A6", -- 0x1508
		x"78",x"86",x"D0",x"90",x"01",x"E8",x"86",x"7A", -- 0x1510
		x"A0",x"00",x"B1",x"79",x"48",x"A9",x"00",x"91", -- 0x1518
		x"79",x"20",x"CE",x"00",x"20",x"31",x"DA",x"68", -- 0x1520
		x"A0",x"00",x"91",x"79",x"A6",x"C6",x"A4",x"C7", -- 0x1528
		x"86",x"CF",x"84",x"D0",x"60",x"20",x"82",x"CB", -- 0x1530
		x"20",x"41",x"D5",x"20",x"DC",x"CC",x"4C",x"E7", -- 0x1538
		x"D4",x"A5",x"BB",x"30",x"9C",x"A5",x"B6",x"C9", -- 0x1540
		x"91",x"B0",x"96",x"20",x"D9",x"D9",x"A5",x"B9", -- 0x1548
		x"A4",x"BA",x"84",x"0E",x"85",x"0F",x"60",x"20", -- 0x1550
		x"41",x"D5",x"A0",x"00",x"B1",x"0E",x"A8",x"4C", -- 0x1558
		x"EF",x"D0",x"20",x"35",x"D5",x"8A",x"A0",x"00", -- 0x1560
		x"91",x"0E",x"60",x"20",x"35",x"D5",x"86",x"9E", -- 0x1568
		x"A2",x"00",x"20",x"CE",x"00",x"F0",x"03",x"20", -- 0x1570
		x"3B",x"D5",x"86",x"9F",x"A0",x"00",x"B1",x"0E", -- 0x1578
		x"45",x"9F",x"25",x"9E",x"F0",x"F8",x"60",x"A9", -- 0x1580
		x"4B",x"A0",x"DC",x"4C",x"A5",x"D5",x"20",x"CA", -- 0x1588
		x"D7",x"A5",x"BB",x"49",x"FF",x"85",x"BB",x"45", -- 0x1590
		x"C3",x"85",x"C4",x"A5",x"B6",x"4C",x"A8",x"D5", -- 0x1598
		x"20",x"D7",x"D6",x"90",x"3C",x"20",x"CA",x"D7", -- 0x15A0
		x"D0",x"03",x"4C",x"3A",x"D9",x"A6",x"C5",x"86", -- 0x15A8
		x"AB",x"A2",x"BE",x"A5",x"BE",x"A8",x"F0",x"CE", -- 0x15B0
		x"38",x"E5",x"B6",x"F0",x"24",x"90",x"12",x"84", -- 0x15B8
		x"B6",x"A4",x"C3",x"84",x"BB",x"49",x"FF",x"69", -- 0x15C0
		x"00",x"A0",x"00",x"84",x"AB",x"A2",x"B6",x"D0", -- 0x15C8
		x"04",x"A0",x"00",x"84",x"C5",x"C9",x"F9",x"30", -- 0x15D0
		x"C7",x"A8",x"A5",x"C5",x"56",x"01",x"20",x"EE", -- 0x15D8
		x"D6",x"24",x"C4",x"10",x"57",x"A0",x"B6",x"E0", -- 0x15E0
		x"BE",x"F0",x"02",x"A0",x"BE",x"38",x"49",x"FF", -- 0x15E8
		x"65",x"AB",x"85",x"C5",x"B9",x"04",x"00",x"F5", -- 0x15F0
		x"04",x"85",x"BA",x"B9",x"03",x"00",x"F5",x"03", -- 0x15F8
		x"85",x"B9",x"B9",x"02",x"00",x"F5",x"02",x"85", -- 0x1600
		x"B8",x"B9",x"01",x"00",x"F5",x"01",x"85",x"B7", -- 0x1608
		x"B0",x"03",x"20",x"85",x"D6",x"A0",x"00",x"98", -- 0x1610
		x"18",x"A6",x"B7",x"D0",x"4A",x"A6",x"B8",x"86", -- 0x1618
		x"B7",x"A6",x"B9",x"86",x"B8",x"A6",x"BA",x"86", -- 0x1620
		x"B9",x"A6",x"C5",x"86",x"BA",x"84",x"C5",x"69", -- 0x1628
		x"08",x"C9",x"20",x"D0",x"E4",x"A9",x"00",x"85", -- 0x1630
		x"B6",x"85",x"BB",x"60",x"65",x"AB",x"85",x"C5", -- 0x1638
		x"A5",x"BA",x"65",x"C2",x"85",x"BA",x"A5",x"B9", -- 0x1640
		x"65",x"C1",x"85",x"B9",x"A5",x"B8",x"65",x"C0", -- 0x1648
		x"85",x"B8",x"A5",x"B7",x"65",x"BF",x"85",x"B7", -- 0x1650
		x"4C",x"74",x"D6",x"69",x"01",x"06",x"C5",x"26", -- 0x1658
		x"BA",x"26",x"B9",x"26",x"B8",x"26",x"B7",x"10", -- 0x1660
		x"F2",x"38",x"E5",x"B6",x"B0",x"C7",x"49",x"FF", -- 0x1668
		x"69",x"01",x"85",x"B6",x"90",x"0E",x"E6",x"B6", -- 0x1670
		x"F0",x"42",x"66",x"B7",x"66",x"B8",x"66",x"B9", -- 0x1678
		x"66",x"BA",x"66",x"C5",x"60",x"A5",x"BB",x"49", -- 0x1680
		x"FF",x"85",x"BB",x"A5",x"B7",x"49",x"FF",x"85", -- 0x1688
		x"B7",x"A5",x"B8",x"49",x"FF",x"85",x"B8",x"A5", -- 0x1690
		x"B9",x"49",x"FF",x"85",x"B9",x"A5",x"BA",x"49", -- 0x1698
		x"FF",x"85",x"BA",x"A5",x"C5",x"49",x"FF",x"85", -- 0x16A0
		x"C5",x"E6",x"C5",x"D0",x"0E",x"E6",x"BA",x"D0", -- 0x16A8
		x"0A",x"E6",x"B9",x"D0",x"06",x"E6",x"B8",x"D0", -- 0x16B0
		x"02",x"E6",x"B7",x"60",x"A2",x"45",x"4C",x"20", -- 0x16B8
		x"C3",x"A2",x"7A",x"B4",x"04",x"84",x"C5",x"B4", -- 0x16C0
		x"03",x"94",x"04",x"B4",x"02",x"94",x"03",x"B4", -- 0x16C8
		x"01",x"94",x"02",x"A4",x"BD",x"94",x"01",x"69", -- 0x16D0
		x"08",x"30",x"E8",x"F0",x"E6",x"E9",x"08",x"A8", -- 0x16D8
		x"A5",x"C5",x"B0",x"14",x"16",x"01",x"90",x"02", -- 0x16E0
		x"F6",x"01",x"76",x"01",x"76",x"01",x"76",x"02", -- 0x16E8
		x"76",x"03",x"76",x"04",x"6A",x"C8",x"D0",x"EC", -- 0x16F0
		x"18",x"60",x"81",x"00",x"00",x"00",x"00",x"03", -- 0x16F8
		x"7F",x"5E",x"56",x"CB",x"79",x"80",x"13",x"9B", -- 0x1700
		x"0B",x"64",x"80",x"76",x"38",x"93",x"16",x"82", -- 0x1708
		x"38",x"AA",x"3B",x"20",x"80",x"35",x"04",x"F3", -- 0x1710
		x"34",x"81",x"35",x"04",x"F3",x"34",x"80",x"80", -- 0x1718
		x"00",x"00",x"00",x"80",x"31",x"72",x"17",x"F8", -- 0x1720
		x"20",x"69",x"D9",x"F0",x"02",x"10",x"03",x"4C", -- 0x1728
		x"96",x"CF",x"A5",x"B6",x"E9",x"7F",x"48",x"A9", -- 0x1730
		x"80",x"85",x"B6",x"A9",x"14",x"A0",x"D7",x"20", -- 0x1738
		x"A5",x"D5",x"A9",x"19",x"A0",x"D7",x"20",x"4D", -- 0x1740
		x"D8",x"A9",x"FA",x"A0",x"D6",x"20",x"8E",x"D5", -- 0x1748
		x"A9",x"FF",x"A0",x"D6",x"20",x"43",x"DD",x"A9", -- 0x1750
		x"1E",x"A0",x"D7",x"20",x"A5",x"D5",x"68",x"20", -- 0x1758
		x"BC",x"DA",x"A9",x"23",x"A0",x"D7",x"20",x"CA", -- 0x1760
		x"D7",x"D0",x"03",x"4C",x"C9",x"D7",x"20",x"F5", -- 0x1768
		x"D7",x"A9",x"00",x"85",x"7B",x"85",x"7C",x"85", -- 0x1770
		x"7D",x"85",x"7E",x"A5",x"C5",x"20",x"97",x"D7", -- 0x1778
		x"A5",x"BA",x"20",x"97",x"D7",x"A5",x"B9",x"20", -- 0x1780
		x"97",x"D7",x"A5",x"B8",x"20",x"97",x"D7",x"A5", -- 0x1788
		x"B7",x"20",x"9C",x"D7",x"4C",x"CD",x"D8",x"D0", -- 0x1790
		x"03",x"4C",x"C1",x"D6",x"4A",x"09",x"80",x"A8", -- 0x1798
		x"90",x"19",x"18",x"A5",x"7E",x"65",x"C2",x"85", -- 0x17A0
		x"7E",x"A5",x"7D",x"65",x"C1",x"85",x"7D",x"A5", -- 0x17A8
		x"7C",x"65",x"C0",x"85",x"7C",x"A5",x"7B",x"65", -- 0x17B0
		x"BF",x"85",x"7B",x"66",x"7B",x"66",x"7C",x"66", -- 0x17B8
		x"7D",x"66",x"7E",x"66",x"C5",x"98",x"4A",x"D0", -- 0x17C0
		x"D6",x"60",x"85",x"77",x"84",x"78",x"A0",x"04", -- 0x17C8
		x"B1",x"77",x"85",x"C2",x"88",x"B1",x"77",x"85", -- 0x17D0
		x"C1",x"88",x"B1",x"77",x"85",x"C0",x"88",x"B1", -- 0x17D8
		x"77",x"85",x"C3",x"45",x"BB",x"85",x"C4",x"A5", -- 0x17E0
		x"C3",x"09",x"80",x"85",x"BF",x"88",x"B1",x"77", -- 0x17E8
		x"85",x"BE",x"A5",x"B6",x"60",x"A5",x"BE",x"F0", -- 0x17F0
		x"1F",x"18",x"65",x"B6",x"90",x"04",x"30",x"1D", -- 0x17F8
		x"18",x"2C",x"10",x"14",x"69",x"80",x"85",x"B6", -- 0x1800
		x"D0",x"03",x"4C",x"39",x"D6",x"A5",x"C4",x"85", -- 0x1808
		x"BB",x"60",x"A5",x"BB",x"49",x"FF",x"30",x"05", -- 0x1810
		x"68",x"68",x"4C",x"35",x"D6",x"4C",x"BC",x"D6", -- 0x1818
		x"20",x"4A",x"D9",x"AA",x"F0",x"10",x"18",x"69", -- 0x1820
		x"02",x"B0",x"F2",x"A2",x"00",x"86",x"C4",x"20", -- 0x1828
		x"B5",x"D5",x"E6",x"B6",x"F0",x"E7",x"60",x"84", -- 0x1830
		x"20",x"00",x"00",x"00",x"20",x"4A",x"D9",x"A9", -- 0x1838
		x"37",x"A0",x"D8",x"A2",x"00",x"86",x"C4",x"20", -- 0x1840
		x"E0",x"D8",x"4C",x"50",x"D8",x"20",x"CA",x"D7", -- 0x1848
		x"F0",x"76",x"20",x"59",x"D9",x"A9",x"00",x"38", -- 0x1850
		x"E5",x"B6",x"85",x"B6",x"20",x"F5",x"D7",x"E6", -- 0x1858
		x"B6",x"F0",x"BA",x"A2",x"FC",x"A9",x"01",x"A4", -- 0x1860
		x"BF",x"C4",x"B7",x"D0",x"10",x"A4",x"C0",x"C4", -- 0x1868
		x"B8",x"D0",x"0A",x"A4",x"C1",x"C4",x"B9",x"D0", -- 0x1870
		x"04",x"A4",x"C2",x"C4",x"BA",x"08",x"2A",x"90", -- 0x1878
		x"09",x"E8",x"95",x"7E",x"F0",x"32",x"10",x"34", -- 0x1880
		x"A9",x"01",x"28",x"B0",x"0E",x"06",x"C2",x"26", -- 0x1888
		x"C1",x"26",x"C0",x"26",x"BF",x"B0",x"E6",x"30", -- 0x1890
		x"CE",x"10",x"E2",x"A8",x"A5",x"C2",x"E5",x"BA", -- 0x1898
		x"85",x"C2",x"A5",x"C1",x"E5",x"B9",x"85",x"C1", -- 0x18A0
		x"A5",x"C0",x"E5",x"B8",x"85",x"C0",x"A5",x"BF", -- 0x18A8
		x"E5",x"B7",x"85",x"BF",x"98",x"4C",x"8D",x"D8", -- 0x18B0
		x"A9",x"40",x"D0",x"CE",x"0A",x"0A",x"0A",x"0A", -- 0x18B8
		x"0A",x"0A",x"85",x"C5",x"28",x"4C",x"CD",x"D8", -- 0x18C0
		x"A2",x"85",x"4C",x"20",x"C3",x"A5",x"7B",x"85", -- 0x18C8
		x"B7",x"A5",x"7C",x"85",x"B8",x"A5",x"7D",x"85", -- 0x18D0
		x"B9",x"A5",x"7E",x"85",x"BA",x"4C",x"15",x"D6", -- 0x18D8
		x"85",x"77",x"84",x"78",x"A0",x"04",x"B1",x"77", -- 0x18E0
		x"85",x"BA",x"88",x"B1",x"77",x"85",x"B9",x"88", -- 0x18E8
		x"B1",x"77",x"85",x"B8",x"88",x"B1",x"77",x"85", -- 0x18F0
		x"BB",x"09",x"80",x"85",x"B7",x"88",x"B1",x"77", -- 0x18F8
		x"85",x"B6",x"84",x"C5",x"60",x"A2",x"B1",x"2C", -- 0x1900
		x"A2",x"AC",x"A0",x"00",x"F0",x"04",x"A6",x"9E", -- 0x1908
		x"A4",x"9F",x"20",x"59",x"D9",x"86",x"77",x"84", -- 0x1910
		x"78",x"A0",x"04",x"A5",x"BA",x"91",x"77",x"88", -- 0x1918
		x"A5",x"B9",x"91",x"77",x"88",x"A5",x"B8",x"91", -- 0x1920
		x"77",x"88",x"A5",x"BB",x"09",x"7F",x"25",x"B7", -- 0x1928
		x"91",x"77",x"88",x"A5",x"B6",x"91",x"77",x"84", -- 0x1930
		x"C5",x"60",x"A5",x"C3",x"85",x"BB",x"A2",x"05", -- 0x1938
		x"B5",x"BD",x"95",x"B5",x"CA",x"D0",x"F9",x"86", -- 0x1940
		x"C5",x"60",x"20",x"59",x"D9",x"A2",x"06",x"B5", -- 0x1948
		x"B5",x"95",x"BD",x"CA",x"D0",x"F9",x"86",x"C5", -- 0x1950
		x"60",x"A5",x"B6",x"F0",x"FB",x"06",x"C5",x"90", -- 0x1958
		x"F7",x"20",x"AD",x"D6",x"D0",x"F2",x"4C",x"76", -- 0x1960
		x"D6",x"A5",x"B6",x"F0",x"09",x"A5",x"BB",x"2A", -- 0x1968
		x"A9",x"FF",x"B0",x"02",x"A9",x"01",x"60",x"20", -- 0x1970
		x"69",x"D9",x"85",x"B7",x"A9",x"00",x"85",x"B8", -- 0x1978
		x"A2",x"88",x"A5",x"B7",x"49",x"FF",x"2A",x"A9", -- 0x1980
		x"00",x"85",x"BA",x"85",x"B9",x"86",x"B6",x"85", -- 0x1988
		x"C5",x"85",x"BB",x"4C",x"10",x"D6",x"46",x"BB", -- 0x1990
		x"60",x"85",x"79",x"84",x"7A",x"A0",x"00",x"B1", -- 0x1998
		x"79",x"C8",x"AA",x"F0",x"C4",x"B1",x"79",x"45", -- 0x19A0
		x"BB",x"30",x"C2",x"E4",x"B6",x"D0",x"21",x"B1", -- 0x19A8
		x"79",x"09",x"80",x"C5",x"B7",x"D0",x"19",x"C8", -- 0x19B0
		x"B1",x"79",x"C5",x"B8",x"D0",x"12",x"C8",x"B1", -- 0x19B8
		x"79",x"C5",x"B9",x"D0",x"0B",x"C8",x"A9",x"7F", -- 0x19C0
		x"C5",x"C5",x"B1",x"79",x"E5",x"BA",x"F0",x"28", -- 0x19C8
		x"A5",x"BB",x"90",x"02",x"49",x"FF",x"4C",x"6F", -- 0x19D0
		x"D9",x"A5",x"B6",x"F0",x"4A",x"38",x"E9",x"A0", -- 0x19D8
		x"24",x"BB",x"10",x"09",x"AA",x"A9",x"FF",x"85", -- 0x19E0
		x"BD",x"20",x"8B",x"D6",x"8A",x"A2",x"B6",x"C9", -- 0x19E8
		x"F9",x"10",x"06",x"20",x"D7",x"D6",x"84",x"BD", -- 0x19F0
		x"60",x"A8",x"A5",x"BB",x"29",x"80",x"46",x"B7", -- 0x19F8
		x"05",x"B7",x"85",x"B7",x"20",x"EE",x"D6",x"84", -- 0x1A00
		x"BD",x"60",x"A5",x"B6",x"C9",x"A0",x"B0",x"20", -- 0x1A08
		x"20",x"D9",x"D9",x"84",x"C5",x"A5",x"BB",x"84", -- 0x1A10
		x"BB",x"49",x"80",x"2A",x"A9",x"A0",x"85",x"B6", -- 0x1A18
		x"A5",x"BA",x"85",x"60",x"4C",x"10",x"D6",x"85", -- 0x1A20
		x"B7",x"85",x"B8",x"85",x"B9",x"85",x"BA",x"A8", -- 0x1A28
		x"60",x"A0",x"00",x"A2",x"0A",x"94",x"B2",x"CA", -- 0x1A30
		x"10",x"FB",x"90",x"0F",x"C9",x"2D",x"D0",x"04", -- 0x1A38
		x"86",x"BC",x"F0",x"04",x"C9",x"2B",x"D0",x"05", -- 0x1A40
		x"20",x"C8",x"00",x"90",x"5B",x"C9",x"2E",x"F0", -- 0x1A48
		x"2E",x"C9",x"45",x"D0",x"30",x"20",x"C8",x"00", -- 0x1A50
		x"90",x"17",x"C9",x"A4",x"F0",x"0E",x"C9",x"2D", -- 0x1A58
		x"F0",x"0A",x"C9",x"A3",x"F0",x"08",x"C9",x"2B", -- 0x1A60
		x"F0",x"04",x"D0",x"07",x"66",x"B5",x"20",x"C8", -- 0x1A68
		x"00",x"90",x"5C",x"24",x"B5",x"10",x"0E",x"A9", -- 0x1A70
		x"00",x"38",x"E5",x"B3",x"4C",x"87",x"DA",x"66", -- 0x1A78
		x"B4",x"24",x"B4",x"50",x"C3",x"A5",x"B3",x"38", -- 0x1A80
		x"E5",x"B2",x"85",x"B3",x"F0",x"12",x"10",x"09", -- 0x1A88
		x"20",x"3C",x"D8",x"E6",x"B3",x"D0",x"F9",x"F0", -- 0x1A90
		x"07",x"20",x"20",x"D8",x"C6",x"B3",x"D0",x"F9", -- 0x1A98
		x"A5",x"BC",x"30",x"01",x"60",x"4C",x"B7",x"DC", -- 0x1AA0
		x"48",x"24",x"B4",x"10",x"02",x"E6",x"B2",x"20", -- 0x1AA8
		x"20",x"D8",x"68",x"38",x"E9",x"30",x"20",x"BC", -- 0x1AB0
		x"DA",x"4C",x"48",x"DA",x"48",x"20",x"4A",x"D9", -- 0x1AB8
		x"68",x"20",x"7A",x"D9",x"A5",x"C3",x"45",x"BB", -- 0x1AC0
		x"85",x"C4",x"A6",x"B6",x"4C",x"A8",x"D5",x"A5", -- 0x1AC8
		x"B3",x"C9",x"0A",x"90",x"09",x"A9",x"64",x"24", -- 0x1AD0
		x"B5",x"30",x"11",x"4C",x"BC",x"D6",x"0A",x"0A", -- 0x1AD8
		x"18",x"65",x"B3",x"0A",x"18",x"A0",x"00",x"71", -- 0x1AE0
		x"CF",x"38",x"E9",x"30",x"85",x"B3",x"4C",x"6E", -- 0x1AE8
		x"DA",x"9B",x"3E",x"BC",x"1F",x"FD",x"9E",x"6E", -- 0x1AF0
		x"6B",x"27",x"FD",x"9E",x"6E",x"6B",x"28",x"00", -- 0x1AF8
		x"A9",x"5F",x"A0",x"C2",x"20",x"18",x"DB",x"A5", -- 0x1B00
		x"8F",x"A6",x"8E",x"85",x"B7",x"86",x"B8",x"A2", -- 0x1B08
		x"90",x"38",x"20",x"87",x"D9",x"20",x"1B",x"DB", -- 0x1B10
		x"4C",x"78",x"C9",x"A0",x"01",x"A9",x"20",x"24", -- 0x1B18
		x"BB",x"10",x"02",x"A9",x"2D",x"99",x"FF",x"00", -- 0x1B20
		x"85",x"BB",x"84",x"C6",x"C8",x"A9",x"30",x"A6", -- 0x1B28
		x"B6",x"D0",x"03",x"4C",x"3E",x"DC",x"A9",x"00", -- 0x1B30
		x"E0",x"80",x"F0",x"02",x"B0",x"09",x"A9",x"FB", -- 0x1B38
		x"A0",x"DA",x"20",x"66",x"D7",x"A9",x"F7",x"85", -- 0x1B40
		x"B2",x"A9",x"F6",x"A0",x"DA",x"20",x"99",x"D9", -- 0x1B48
		x"F0",x"1E",x"10",x"12",x"A9",x"F1",x"A0",x"DA", -- 0x1B50
		x"20",x"99",x"D9",x"F0",x"02",x"10",x"0E",x"20", -- 0x1B58
		x"20",x"D8",x"C6",x"B2",x"D0",x"EE",x"20",x"3C", -- 0x1B60
		x"D8",x"E6",x"B2",x"D0",x"DC",x"20",x"87",x"D5", -- 0x1B68
		x"20",x"D9",x"D9",x"A2",x"01",x"A5",x"B2",x"18", -- 0x1B70
		x"69",x"0A",x"30",x"09",x"C9",x"0B",x"B0",x"06", -- 0x1B78
		x"69",x"FF",x"AA",x"A9",x"02",x"38",x"E9",x"02", -- 0x1B80
		x"85",x"B3",x"86",x"B2",x"8A",x"F0",x"02",x"10", -- 0x1B88
		x"13",x"A4",x"C6",x"A9",x"2E",x"C8",x"99",x"FF", -- 0x1B90
		x"00",x"8A",x"F0",x"06",x"A9",x"30",x"C8",x"99", -- 0x1B98
		x"FF",x"00",x"84",x"C6",x"A0",x"00",x"A2",x"80", -- 0x1BA0
		x"A5",x"BA",x"18",x"79",x"53",x"DC",x"85",x"BA", -- 0x1BA8
		x"A5",x"B9",x"79",x"52",x"DC",x"85",x"B9",x"A5", -- 0x1BB0
		x"B8",x"79",x"51",x"DC",x"85",x"B8",x"A5",x"B7", -- 0x1BB8
		x"79",x"50",x"DC",x"85",x"B7",x"E8",x"B0",x"04", -- 0x1BC0
		x"10",x"DE",x"30",x"02",x"30",x"DA",x"8A",x"90", -- 0x1BC8
		x"04",x"49",x"FF",x"69",x"0A",x"69",x"2F",x"C8", -- 0x1BD0
		x"C8",x"C8",x"C8",x"84",x"9C",x"A4",x"C6",x"C8", -- 0x1BD8
		x"AA",x"29",x"7F",x"99",x"FF",x"00",x"C6",x"B2", -- 0x1BE0
		x"D0",x"06",x"A9",x"2E",x"C8",x"99",x"FF",x"00", -- 0x1BE8
		x"84",x"C6",x"A4",x"9C",x"8A",x"49",x"FF",x"29", -- 0x1BF0
		x"80",x"AA",x"C0",x"24",x"D0",x"AA",x"A4",x"C6", -- 0x1BF8
		x"B9",x"FF",x"00",x"88",x"C9",x"30",x"F0",x"F8", -- 0x1C00
		x"C9",x"2E",x"F0",x"01",x"C8",x"A9",x"2B",x"A6", -- 0x1C08
		x"B3",x"F0",x"2E",x"10",x"08",x"A9",x"00",x"38", -- 0x1C10
		x"E5",x"B3",x"AA",x"A9",x"2D",x"99",x"01",x"01", -- 0x1C18
		x"A9",x"45",x"99",x"00",x"01",x"8A",x"A2",x"2F", -- 0x1C20
		x"38",x"E8",x"E9",x"0A",x"B0",x"FB",x"69",x"3A", -- 0x1C28
		x"99",x"03",x"01",x"8A",x"99",x"02",x"01",x"A9", -- 0x1C30
		x"00",x"99",x"04",x"01",x"F0",x"08",x"99",x"FF", -- 0x1C38
		x"00",x"A9",x"00",x"99",x"00",x"01",x"A9",x"00", -- 0x1C40
		x"A0",x"01",x"60",x"80",x"00",x"00",x"00",x"00", -- 0x1C48
		x"FA",x"0A",x"1F",x"00",x"00",x"98",x"96",x"80", -- 0x1C50
		x"FF",x"F0",x"BD",x"C0",x"00",x"01",x"86",x"A0", -- 0x1C58
		x"FF",x"FF",x"D8",x"F0",x"00",x"00",x"03",x"E8", -- 0x1C60
		x"FF",x"FF",x"FF",x"9C",x"00",x"00",x"00",x"0A", -- 0x1C68
		x"FF",x"FF",x"FF",x"FF",x"20",x"4A",x"D9",x"A9", -- 0x1C70
		x"4B",x"A0",x"DC",x"20",x"E0",x"D8",x"F0",x"70", -- 0x1C78
		x"A5",x"BE",x"D0",x"03",x"4C",x"37",x"D6",x"A2", -- 0x1C80
		x"A3",x"A0",x"00",x"20",x"12",x"D9",x"A5",x"C3", -- 0x1C88
		x"10",x"0F",x"20",x"0A",x"DA",x"A9",x"A3",x"A0", -- 0x1C90
		x"00",x"20",x"99",x"D9",x"D0",x"03",x"98",x"A4", -- 0x1C98
		x"60",x"20",x"3C",x"D9",x"98",x"48",x"20",x"28", -- 0x1CA0
		x"D7",x"A9",x"A3",x"A0",x"00",x"20",x"66",x"D7", -- 0x1CA8
		x"20",x"F0",x"DC",x"68",x"4A",x"90",x"0A",x"A5", -- 0x1CB0
		x"B6",x"F0",x"06",x"A5",x"BB",x"49",x"FF",x"85", -- 0x1CB8
		x"BB",x"60",x"81",x"38",x"AA",x"3B",x"29",x"07", -- 0x1CC0
		x"71",x"34",x"58",x"3E",x"56",x"74",x"16",x"7E", -- 0x1CC8
		x"B3",x"1B",x"77",x"2F",x"EE",x"E3",x"85",x"7A", -- 0x1CD0
		x"1D",x"84",x"1C",x"2A",x"7C",x"63",x"59",x"58", -- 0x1CD8
		x"0A",x"7E",x"75",x"FD",x"E7",x"C6",x"80",x"31", -- 0x1CE0
		x"72",x"18",x"10",x"81",x"00",x"00",x"00",x"00", -- 0x1CE8
		x"A9",x"C2",x"A0",x"DC",x"20",x"66",x"D7",x"A5", -- 0x1CF0
		x"C5",x"69",x"50",x"90",x"03",x"20",x"61",x"D9", -- 0x1CF8
		x"85",x"AB",x"20",x"4D",x"D9",x"A5",x"B6",x"C9", -- 0x1D00
		x"88",x"90",x"03",x"20",x"12",x"D8",x"20",x"0A", -- 0x1D08
		x"DA",x"A5",x"60",x"18",x"69",x"81",x"F0",x"F3", -- 0x1D10
		x"38",x"E9",x"01",x"48",x"A2",x"05",x"B5",x"BE", -- 0x1D18
		x"B4",x"B6",x"95",x"B6",x"94",x"BE",x"CA",x"10", -- 0x1D20
		x"F5",x"A5",x"AB",x"85",x"C5",x"20",x"91",x"D5", -- 0x1D28
		x"20",x"B7",x"DC",x"A9",x"C7",x"A0",x"DC",x"20", -- 0x1D30
		x"59",x"DD",x"A9",x"00",x"85",x"C4",x"68",x"20", -- 0x1D38
		x"F7",x"D7",x"60",x"85",x"C6",x"84",x"C7",x"20", -- 0x1D40
		x"08",x"D9",x"A9",x"AC",x"20",x"66",x"D7",x"20", -- 0x1D48
		x"5D",x"DD",x"A9",x"AC",x"A0",x"00",x"4C",x"66", -- 0x1D50
		x"D7",x"85",x"C6",x"84",x"C7",x"20",x"05",x"D9", -- 0x1D58
		x"B1",x"C6",x"85",x"BC",x"A4",x"C6",x"C8",x"98", -- 0x1D60
		x"D0",x"02",x"E6",x"C7",x"85",x"C6",x"A4",x"C7", -- 0x1D68
		x"20",x"66",x"D7",x"A5",x"C6",x"A4",x"C7",x"18", -- 0x1D70
		x"69",x"05",x"90",x"01",x"C8",x"85",x"C6",x"84", -- 0x1D78
		x"C7",x"20",x"A5",x"D5",x"A9",x"B1",x"A0",x"00", -- 0x1D80
		x"C6",x"BC",x"D0",x"E4",x"60",x"98",x"35",x"44", -- 0x1D88
		x"7A",x"68",x"28",x"B1",x"46",x"20",x"69",x"D9", -- 0x1D90
		x"AA",x"30",x"18",x"A9",x"E0",x"A0",x"00",x"20", -- 0x1D98
		x"E0",x"D8",x"8A",x"F0",x"E7",x"A9",x"8D",x"A0", -- 0x1DA0
		x"DD",x"20",x"66",x"D7",x"A9",x"91",x"A0",x"DD", -- 0x1DA8
		x"20",x"A5",x"D5",x"A6",x"BA",x"A5",x"B7",x"85", -- 0x1DB0
		x"BA",x"86",x"B7",x"A9",x"00",x"85",x"BB",x"A5", -- 0x1DB8
		x"B6",x"85",x"C5",x"A9",x"80",x"85",x"B6",x"20", -- 0x1DC0
		x"15",x"D6",x"A2",x"E0",x"A0",x"00",x"4C",x"12", -- 0x1DC8
		x"D9",x"A9",x"4D",x"A0",x"DE",x"20",x"A5",x"D5", -- 0x1DD0
		x"20",x"4A",x"D9",x"A9",x"52",x"A0",x"DE",x"A6", -- 0x1DD8
		x"C3",x"20",x"45",x"D8",x"20",x"4A",x"D9",x"20", -- 0x1DE0
		x"0A",x"DA",x"A9",x"00",x"85",x"C4",x"20",x"91", -- 0x1DE8
		x"D5",x"A9",x"57",x"A0",x"DE",x"20",x"8E",x"D5", -- 0x1DF0
		x"A5",x"BB",x"48",x"10",x"0D",x"20",x"87",x"D5", -- 0x1DF8
		x"A5",x"BB",x"30",x"09",x"A5",x"69",x"49",x"FF", -- 0x1E00
		x"85",x"69",x"20",x"B7",x"DC",x"A9",x"57",x"A0", -- 0x1E08
		x"DE",x"20",x"A5",x"D5",x"68",x"10",x"03",x"20", -- 0x1E10
		x"B7",x"DC",x"A9",x"5C",x"A0",x"DE",x"4C",x"43", -- 0x1E18
		x"DD",x"20",x"08",x"D9",x"A9",x"00",x"85",x"69", -- 0x1E20
		x"20",x"D8",x"DD",x"A2",x"A3",x"A0",x"00",x"20", -- 0x1E28
		x"CE",x"DD",x"A9",x"AC",x"A0",x"00",x"20",x"E0", -- 0x1E30
		x"D8",x"A9",x"00",x"85",x"BB",x"A5",x"69",x"20", -- 0x1E38
		x"49",x"DE",x"A9",x"A3",x"A0",x"00",x"4C",x"4D", -- 0x1E40
		x"D8",x"48",x"4C",x"0A",x"DE",x"81",x"49",x"0F", -- 0x1E48
		x"DA",x"A2",x"83",x"49",x"0F",x"DA",x"A2",x"7F", -- 0x1E50
		x"00",x"00",x"00",x"00",x"05",x"84",x"E6",x"1A", -- 0x1E58
		x"2D",x"1B",x"86",x"28",x"07",x"FB",x"F8",x"87", -- 0x1E60
		x"99",x"68",x"89",x"01",x"87",x"23",x"35",x"DF", -- 0x1E68
		x"E1",x"86",x"A5",x"5D",x"E7",x"28",x"83",x"49", -- 0x1E70
		x"0F",x"DA",x"A2",x"A1",x"54",x"46",x"8F",x"13", -- 0x1E78
		x"8F",x"52",x"43",x"89",x"CD",x"A5",x"BB",x"48", -- 0x1E80
		x"10",x"03",x"20",x"B7",x"DC",x"A5",x"B6",x"48", -- 0x1E88
		x"C9",x"81",x"90",x"07",x"A9",x"FA",x"A0",x"D6", -- 0x1E90
		x"20",x"4D",x"D8",x"A9",x"B5",x"A0",x"DE",x"20", -- 0x1E98
		x"43",x"DD",x"68",x"C9",x"81",x"90",x"07",x"A9", -- 0x1EA0
		x"4D",x"A0",x"DE",x"20",x"8E",x"D5",x"68",x"10", -- 0x1EA8
		x"03",x"4C",x"B7",x"DC",x"60",x"0B",x"76",x"B3", -- 0x1EB0
		x"83",x"BD",x"D3",x"79",x"1E",x"F4",x"A6",x"F5", -- 0x1EB8
		x"7B",x"83",x"FC",x"B0",x"10",x"7C",x"0C",x"1F", -- 0x1EC0
		x"67",x"CA",x"7C",x"DE",x"53",x"CB",x"C1",x"7D", -- 0x1EC8
		x"14",x"64",x"70",x"4C",x"7D",x"B7",x"EA",x"51", -- 0x1ED0
		x"7A",x"7D",x"63",x"30",x"88",x"7E",x"7E",x"92", -- 0x1ED8
		x"44",x"99",x"3A",x"7E",x"4C",x"CC",x"91",x"C7", -- 0x1EE0
		x"7F",x"AA",x"AA",x"AA",x"13",x"81",x"00",x"00", -- 0x1EE8
		x"00",x"00",x"E6",x"CF",x"D0",x"02",x"E6",x"D0", -- 0x1EF0
		x"AD",x"60",x"EA",x"C9",x"3A",x"B0",x"0A",x"C9", -- 0x1EF8
		x"20",x"F0",x"EF",x"38",x"E9",x"30",x"38",x"E9", -- 0x1F00
		x"D0",x"60",x"80",x"4F",x"C7",x"52",x"58",x"A9", -- 0x1F08
		x"3E",x"A0",x"E0",x"20",x"78",x"C9",x"A2",x"FF", -- 0x1F10
		x"86",x"8F",x"9A",x"A9",x"16",x"A0",x"DF",x"85", -- 0x1F18
		x"01",x"84",x"02",x"85",x"04",x"84",x"05",x"A9", -- 0x1F20
		x"0D",x"A0",x"CF",x"85",x"06",x"84",x"07",x"A9", -- 0x1F28
		x"E0",x"A0",x"D0",x"85",x"08",x"84",x"09",x"A9", -- 0x1F30
		x"4C",x"85",x"00",x"85",x"03",x"85",x"A9",x"85", -- 0x1F38
		x"00",x"A9",x"96",x"A0",x"CF",x"85",x"01",x"84", -- 0x1F40
		x"02",x"A9",x"28",x"85",x"0C",x"A9",x"1E",x"85", -- 0x1F48
		x"0D",x"A2",x"1C",x"BD",x"F1",x"DE",x"95",x"C7", -- 0x1F50
		x"CA",x"D0",x"F8",x"A9",x"03",x"85",x"A8",x"8A", -- 0x1F58
		x"85",x"BD",x"85",x"6D",x"48",x"85",x"6A",x"A9", -- 0x1F60
		x"03",x"85",x"A8",x"20",x"32",x"C9",x"A2",x"6E", -- 0x1F68
		x"86",x"6B",x"A9",x"5E",x"A0",x"E0",x"20",x"78", -- 0x1F70
		x"C9",x"20",x"01",x"CA",x"86",x"CF",x"84",x"D0", -- 0x1F78
		x"20",x"C8",x"00",x"C9",x"41",x"F0",x"88",x"A8", -- 0x1F80
		x"D0",x"25",x"A9",x"00",x"A0",x"04",x"85",x"80", -- 0x1F88
		x"84",x"81",x"85",x"0E",x"84",x"0F",x"A0",x"00", -- 0x1F90
		x"E6",x"0E",x"D0",x"02",x"E6",x"0F",x"A9",x"55", -- 0x1F98
		x"91",x"0E",x"D1",x"0E",x"D0",x"15",x"0A",x"91", -- 0x1FA0
		x"0E",x"D1",x"0E",x"D0",x"0E",x"F0",x"E9",x"20", -- 0x1FA8
		x"CE",x"00",x"20",x"2B",x"C8",x"A8",x"F0",x"03", -- 0x1FB0
		x"4C",x"E7",x"CC",x"A5",x"0E",x"A4",x"0F",x"85", -- 0x1FB8
		x"8C",x"84",x"8D",x"85",x"88",x"84",x"89",x"A9", -- 0x1FC0
		x"6A",x"A0",x"E0",x"20",x"78",x"C9",x"20",x"01", -- 0x1FC8
		x"CA",x"86",x"CF",x"84",x"D0",x"20",x"C8",x"00", -- 0x1FD0
		x"A8",x"F0",x"1C",x"20",x"2B",x"C8",x"A5",x"0F", -- 0x1FD8
		x"D0",x"E5",x"A5",x"0E",x"C9",x"10",x"90",x"DF", -- 0x1FE0
		x"85",x"0C",x"E9",x"0E",x"B0",x"FC",x"49",x"FF", -- 0x1FE8
		x"E9",x"0C",x"18",x"65",x"0C",x"85",x"0D",x"A2", -- 0x1FF0
		x"00",x"A0",x"04",x"86",x"80",x"84",x"81",x"A0", -- 0x1FF8
		x"00",x"98",x"91",x"80",x"E6",x"80",x"D0",x"02", -- 0x2000
		x"E6",x"81",x"A5",x"80",x"A4",x"81",x"20",x"F1", -- 0x2008
		x"C2",x"20",x"32",x"C9",x"A5",x"8C",x"38",x"E5", -- 0x2010
		x"80",x"AA",x"A5",x"8D",x"E5",x"81",x"20",x"0B", -- 0x2018
		x"DB",x"A9",x"79",x"A0",x"E0",x"20",x"78",x"C9", -- 0x2020
		x"20",x"25",x"C5",x"A9",x"78",x"A0",x"C9",x"85", -- 0x2028
		x"04",x"84",x"05",x"A9",x"47",x"A0",x"C3",x"85", -- 0x2030
		x"01",x"84",x"02",x"6C",x"01",x"00",x"0D",x"0A", -- 0x2038
		x"0C",x"57",x"52",x"49",x"54",x"54",x"45",x"4E", -- 0x2040
		x"20",x"42",x"59",x"20",x"57",x"45",x"49",x"4C", -- 0x2048
		x"41",x"4E",x"44",x"20",x"26",x"20",x"47",x"41", -- 0x2050
		x"54",x"45",x"53",x"0D",x"0A",x"00",x"4D",x"45", -- 0x2058
		x"4D",x"4F",x"52",x"59",x"20",x"53",x"49",x"5A", -- 0x2060
		x"45",x"00",x"54",x"45",x"52",x"4D",x"49",x"4E", -- 0x2068
		x"41",x"4C",x"20",x"57",x"49",x"44",x"54",x"48", -- 0x2070
		x"00",x"20",x"42",x"59",x"54",x"45",x"53",x"20", -- 0x2078
		x"46",x"52",x"45",x"45",x"0D",x"0A",x"0D",x"0A", -- 0x2080
		x"0D",x"0A",x"43",x"4F",x"50",x"59",x"52",x"49", -- 0x2088
		x"47",x"48",x"54",x"20",x"31",x"39",x"37",x"37", -- 0x2090
		x"20",x"42",x"59",x"20",x"4D",x"49",x"43",x"52", -- 0x2098
		x"4F",x"53",x"4F",x"46",x"54",x"20",x"43",x"4F", -- 0x20A0
		x"2E",x"0D",x"0A",x"00",x"00",x"00",x"00",x"00", -- 0x20A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2100
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2108
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2110
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2118
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2120
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2128
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2130
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2138
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2140
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2148
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2150
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2158
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2160
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2168
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2170
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2178
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2180
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2188
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2190
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2198
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x21A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x21A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x21B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x21B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x21C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x21C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x21D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x21D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x21E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x21E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x21F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x21F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2200
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2208
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2210
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2218
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2220
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2228
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2230
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2238
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2240
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2248
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2250
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2258
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2260
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2268
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2270
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2278
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2280
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2288
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2290
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2298
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x22A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x22A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x22B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x22B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x22C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x22C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x22D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x22D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x22E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x22E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x22F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x22F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2300
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2308
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2310
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2318
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2320
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2328
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2330
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2338
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2340
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2348
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2350
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2358
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2360
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2368
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2370
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2378
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2380
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2388
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2390
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2398
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x23A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x23A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x23B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x23B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x23C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x23C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x23D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x23D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x23E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x23E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x23F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x23F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2400
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2408
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2410
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2418
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2420
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2428
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2430
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2438
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2440
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2448
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2450
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2458
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2460
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2468
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2470
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2478
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2480
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2488
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2490
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2498
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x24F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2500
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2508
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2510
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2518
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2520
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2528
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2530
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2538
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2540
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2548
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2550
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2558
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2560
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2568
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2570
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2578
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2580
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2588
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2590
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2598
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x25F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2600
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2608
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2610
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2618
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2620
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2628
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2630
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2638
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2640
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2648
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2650
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2658
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2660
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2668
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2670
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2678
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2680
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2688
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2690
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2698
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x26A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x26A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x26B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x26B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x26C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x26C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x26D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x26D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x26E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x26E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x26F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x26F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2700
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2708
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2710
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2718
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2720
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2728
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2730
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2738
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2740
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2748
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2750
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2758
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2760
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2768
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2770
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2778
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2780
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2788
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2790
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2798
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x27A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x27A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x27B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x27B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x27C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x27C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x27D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x27D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x27E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x27E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x27F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x27F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2800
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2808
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2810
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2818
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2820
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2828
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2830
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2838
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2840
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2848
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2850
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2858
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2860
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2868
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2870
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2878
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2880
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2888
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2890
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2898
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2900
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2908
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2910
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2918
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2920
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2928
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2930
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2938
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2940
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2948
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2950
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2958
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2960
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2968
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2970
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2978
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2980
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2988
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2990
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2998
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2ED0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2ED8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3000
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3008
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3010
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3018
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3020
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3028
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3030
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3038
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3040
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3048
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3050
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3058
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3060
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3068
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3070
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3078
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3080
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3088
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3090
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3098
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3100
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3108
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3110
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3118
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3120
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3128
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3130
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3138
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3140
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3148
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3150
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3158
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3160
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3168
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3170
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3178
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3180
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3188
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3190
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3198
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3200
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3208
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3210
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3218
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3220
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3228
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3230
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3238
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3240
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3248
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3250
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3258
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3260
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3268
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3270
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3278
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3280
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3288
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3290
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3298
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3300
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3308
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3310
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3318
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3320
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3328
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3330
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3338
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3340
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3348
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3350
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3358
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3360
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3368
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3370
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3378
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3380
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3388
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3390
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3398
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3400
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3408
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3410
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3418
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3420
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3428
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3430
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3438
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3440
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3448
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3450
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3458
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3460
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3468
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3470
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3478
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3480
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3488
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3490
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3498
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3500
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3508
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3510
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3518
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3520
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3528
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3530
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3538
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3540
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3548
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3550
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3558
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3560
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3568
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3570
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3578
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3580
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3588
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3590
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3598
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3600
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3608
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3610
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3618
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3620
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3628
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3630
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3638
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3640
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3648
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3650
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3658
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3660
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3668
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3670
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3678
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3680
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3688
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3690
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3698
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3700
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3708
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3710
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3718
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3720
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3728
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3730
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3738
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3740
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3748
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3750
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3758
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3760
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3768
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3770
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3778
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3780
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3788
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3790
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3798
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3800
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3808
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3810
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3818
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3820
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3828
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3830
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3838
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3840
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3848
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3850
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3858
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3860
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3868
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3870
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3878
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3880
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3888
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3890
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3898
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3900
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3908
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3910
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3918
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3920
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3928
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3930
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3938
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3940
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3948
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3950
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3958
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3960
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3968
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3970
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3978
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3980
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3988
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3990
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3998
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DF8
		x"A0",x"7F",x"C9",x"08",x"F0",x"18",x"C9",x"1B", -- 0x3E00
		x"F0",x"03",x"C8",x"10",x"14",x"A9",x"5C",x"20", -- 0x3E08
		x"FC",x"FE",x"A9",x"0D",x"20",x"FC",x"FE",x"A9", -- 0x3E10
		x"0A",x"20",x"FC",x"FE",x"A0",x"01",x"88",x"30", -- 0x3E18
		x"F1",x"AD",x"E1",x"FC",x"29",x"01",x"F0",x"06", -- 0x3E20
		x"AD",x"E0",x"FC",x"4C",x"38",x"FE",x"AD",x"E3", -- 0x3E28
		x"FC",x"29",x"01",x"F0",x"EC",x"AD",x"E2",x"FC", -- 0x3E30
		x"99",x"00",x"02",x"20",x"FC",x"FE",x"C9",x"0D", -- 0x3E38
		x"D0",x"C0",x"A0",x"FF",x"A9",x"00",x"AA",x"0A", -- 0x3E40
		x"0A",x"85",x"2B",x"C8",x"B9",x"00",x"02",x"C9", -- 0x3E48
		x"0D",x"F0",x"BF",x"C9",x"2E",x"90",x"F4",x"F0", -- 0x3E50
		x"EE",x"C9",x"3A",x"F0",x"EB",x"C9",x"52",x"F0", -- 0x3E58
		x"3B",x"86",x"28",x"86",x"29",x"84",x"2A",x"B9", -- 0x3E60
		x"00",x"02",x"49",x"30",x"C9",x"0A",x"90",x"06", -- 0x3E68
		x"69",x"88",x"C9",x"FA",x"90",x"11",x"0A",x"0A", -- 0x3E70
		x"0A",x"0A",x"A2",x"04",x"0A",x"26",x"28",x"26", -- 0x3E78
		x"29",x"CA",x"D0",x"F8",x"C8",x"D0",x"E0",x"C4", -- 0x3E80
		x"2A",x"F0",x"82",x"24",x"2B",x"50",x"10",x"A5", -- 0x3E88
		x"28",x"81",x"26",x"E6",x"26",x"D0",x"B5",x"E6", -- 0x3E90
		x"27",x"4C",x"4C",x"FE",x"6C",x"24",x"00",x"30", -- 0x3E98
		x"30",x"A2",x"02",x"B5",x"27",x"95",x"25",x"95", -- 0x3EA0
		x"23",x"CA",x"D0",x"F7",x"D0",x"19",x"A9",x"0D", -- 0x3EA8
		x"20",x"FC",x"FE",x"A9",x"0A",x"20",x"FC",x"FE", -- 0x3EB0
		x"A5",x"25",x"20",x"E9",x"FE",x"A5",x"24",x"20", -- 0x3EB8
		x"E9",x"FE",x"A9",x"3A",x"20",x"FC",x"FE",x"A9", -- 0x3EC0
		x"20",x"20",x"FC",x"FE",x"A1",x"24",x"20",x"E9", -- 0x3EC8
		x"FE",x"86",x"2B",x"A5",x"24",x"C5",x"28",x"A5", -- 0x3ED0
		x"25",x"E5",x"29",x"B0",x"BC",x"E6",x"24",x"D0", -- 0x3ED8
		x"02",x"E6",x"25",x"A5",x"24",x"29",x"07",x"10", -- 0x3EE0
		x"C3",x"48",x"4A",x"4A",x"4A",x"4A",x"20",x"F2", -- 0x3EE8
		x"FE",x"68",x"29",x"0F",x"09",x"30",x"C9",x"3A", -- 0x3EF0
		x"90",x"02",x"69",x"06",x"48",x"8D",x"E0",x"FF", -- 0x3EF8
		x"A9",x"FF",x"3A",x"D0",x"FD",x"68",x"60",x"AD", -- 0x3F00
		x"E1",x"FC",x"29",x"01",x"F0",x"08",x"AD",x"E0", -- 0x3F08
		x"FC",x"20",x"FC",x"FE",x"38",x"60",x"AD",x"E3", -- 0x3F10
		x"FC",x"29",x"01",x"F0",x"08",x"AD",x"E2",x"FC", -- 0x3F18
		x"20",x"FC",x"FE",x"38",x"60",x"18",x"60",x"60", -- 0x3F20
		x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FF0
		x"00",x"00",x"00",x"0F",x"00",x"FE",x"00",x"00"  -- 0x3FF8
	);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			data <= rom(to_integer(unsigned(addr)));
		end if;
	end process;
end rtl;
